module wallace_26x26 (
    input  [25:0] a,
    input  [25:0] b,
    output [51:0] p
);

    wire [25:0] pp[25:0];
    genvar i,j;
    generate
        for (i = 0; i < 26; i = i + 1) begin
            for (j = 0; j < 26; j = j + 1) begin
                assign pp[i][j] = a[j] & b[i];
            end
        end
    endgenerate

    wire s_0_2_0, c_0_2_0;
    csa u_csa_0_2_0(pp[2][0],pp[1][1],pp[0][2],s_0_2_0,c_0_2_0);
    wire s_0_3_1, c_0_3_1;
    csa u_csa_0_3_1(pp[3][0],pp[2][1],pp[1][2],s_0_3_1,c_0_3_1);
    wire s_0_4_1, c_0_4_1;
    csa u_csa_0_4_1(pp[4][0],pp[3][1],pp[2][2],s_0_4_1,c_0_4_1);
    wire s_0_5_1, c_0_5_1;
    csa u_csa_0_5_1(pp[5][0],pp[4][1],pp[3][2],s_0_5_1,c_0_5_1);
    wire s_0_5_2, c_0_5_2;
    csa u_csa_0_5_2(pp[2][3],pp[1][4],pp[0][5],s_0_5_2,c_0_5_2);
    wire s_0_6_2, c_0_6_2;
    csa u_csa_0_6_2(pp[6][0],pp[5][1],pp[4][2],s_0_6_2,c_0_6_2);
    wire s_0_6_3, c_0_6_3;
    csa u_csa_0_6_3(pp[3][3],pp[2][4],pp[1][5],s_0_6_3,c_0_6_3);
    wire s_0_7_2, c_0_7_2;
    csa u_csa_0_7_2(pp[7][0],pp[6][1],pp[5][2],s_0_7_2,c_0_7_2);
    wire s_0_7_3, c_0_7_3;
    csa u_csa_0_7_3(pp[4][3],pp[3][4],pp[2][5],s_0_7_3,c_0_7_3);
    wire s_0_8_2, c_0_8_2;
    csa u_csa_0_8_2(pp[8][0],pp[7][1],pp[6][2],s_0_8_2,c_0_8_2);
    wire s_0_8_3, c_0_8_3;
    csa u_csa_0_8_3(pp[5][3],pp[4][4],pp[3][5],s_0_8_3,c_0_8_3);
    wire s_0_8_4, c_0_8_4;
    csa u_csa_0_8_4(pp[2][6],pp[1][7],pp[0][8],s_0_8_4,c_0_8_4);
    wire s_0_9_3, c_0_9_3;
    csa u_csa_0_9_3(pp[9][0],pp[8][1],pp[7][2],s_0_9_3,c_0_9_3);
    wire s_0_9_4, c_0_9_4;
    csa u_csa_0_9_4(pp[6][3],pp[5][4],pp[4][5],s_0_9_4,c_0_9_4);
    wire s_0_9_5, c_0_9_5;
    csa u_csa_0_9_5(pp[3][6],pp[2][7],pp[1][8],s_0_9_5,c_0_9_5);
    wire s_0_10_3, c_0_10_3;
    csa u_csa_0_10_3(pp[10][0],pp[9][1],pp[8][2],s_0_10_3,c_0_10_3);
    wire s_0_10_4, c_0_10_4;
    csa u_csa_0_10_4(pp[7][3],pp[6][4],pp[5][5],s_0_10_4,c_0_10_4);
    wire s_0_10_5, c_0_10_5;
    csa u_csa_0_10_5(pp[4][6],pp[3][7],pp[2][8],s_0_10_5,c_0_10_5);
    wire s_0_11_3, c_0_11_3;
    csa u_csa_0_11_3(pp[11][0],pp[10][1],pp[9][2],s_0_11_3,c_0_11_3);
    wire s_0_11_4, c_0_11_4;
    csa u_csa_0_11_4(pp[8][3],pp[7][4],pp[6][5],s_0_11_4,c_0_11_4);
    wire s_0_11_5, c_0_11_5;
    csa u_csa_0_11_5(pp[5][6],pp[4][7],pp[3][8],s_0_11_5,c_0_11_5);
    wire s_0_11_6, c_0_11_6;
    csa u_csa_0_11_6(pp[2][9],pp[1][10],pp[0][11],s_0_11_6,c_0_11_6);
    wire s_0_12_4, c_0_12_4;
    csa u_csa_0_12_4(pp[12][0],pp[11][1],pp[10][2],s_0_12_4,c_0_12_4);
    wire s_0_12_5, c_0_12_5;
    csa u_csa_0_12_5(pp[9][3],pp[8][4],pp[7][5],s_0_12_5,c_0_12_5);
    wire s_0_12_6, c_0_12_6;
    csa u_csa_0_12_6(pp[6][6],pp[5][7],pp[4][8],s_0_12_6,c_0_12_6);
    wire s_0_12_7, c_0_12_7;
    csa u_csa_0_12_7(pp[3][9],pp[2][10],pp[1][11],s_0_12_7,c_0_12_7);
    wire s_0_13_4, c_0_13_4;
    csa u_csa_0_13_4(pp[13][0],pp[12][1],pp[11][2],s_0_13_4,c_0_13_4);
    wire s_0_13_5, c_0_13_5;
    csa u_csa_0_13_5(pp[10][3],pp[9][4],pp[8][5],s_0_13_5,c_0_13_5);
    wire s_0_13_6, c_0_13_6;
    csa u_csa_0_13_6(pp[7][6],pp[6][7],pp[5][8],s_0_13_6,c_0_13_6);
    wire s_0_13_7, c_0_13_7;
    csa u_csa_0_13_7(pp[4][9],pp[3][10],pp[2][11],s_0_13_7,c_0_13_7);
    wire s_0_14_4, c_0_14_4;
    csa u_csa_0_14_4(pp[14][0],pp[13][1],pp[12][2],s_0_14_4,c_0_14_4);
    wire s_0_14_5, c_0_14_5;
    csa u_csa_0_14_5(pp[11][3],pp[10][4],pp[9][5],s_0_14_5,c_0_14_5);
    wire s_0_14_6, c_0_14_6;
    csa u_csa_0_14_6(pp[8][6],pp[7][7],pp[6][8],s_0_14_6,c_0_14_6);
    wire s_0_14_7, c_0_14_7;
    csa u_csa_0_14_7(pp[5][9],pp[4][10],pp[3][11],s_0_14_7,c_0_14_7);
    wire s_0_14_8, c_0_14_8;
    csa u_csa_0_14_8(pp[2][12],pp[1][13],pp[0][14],s_0_14_8,c_0_14_8);
    wire s_0_15_5, c_0_15_5;
    csa u_csa_0_15_5(pp[15][0],pp[14][1],pp[13][2],s_0_15_5,c_0_15_5);
    wire s_0_15_6, c_0_15_6;
    csa u_csa_0_15_6(pp[12][3],pp[11][4],pp[10][5],s_0_15_6,c_0_15_6);
    wire s_0_15_7, c_0_15_7;
    csa u_csa_0_15_7(pp[9][6],pp[8][7],pp[7][8],s_0_15_7,c_0_15_7);
    wire s_0_15_8, c_0_15_8;
    csa u_csa_0_15_8(pp[6][9],pp[5][10],pp[4][11],s_0_15_8,c_0_15_8);
    wire s_0_15_9, c_0_15_9;
    csa u_csa_0_15_9(pp[3][12],pp[2][13],pp[1][14],s_0_15_9,c_0_15_9);
    wire s_0_16_5, c_0_16_5;
    csa u_csa_0_16_5(pp[16][0],pp[15][1],pp[14][2],s_0_16_5,c_0_16_5);
    wire s_0_16_6, c_0_16_6;
    csa u_csa_0_16_6(pp[13][3],pp[12][4],pp[11][5],s_0_16_6,c_0_16_6);
    wire s_0_16_7, c_0_16_7;
    csa u_csa_0_16_7(pp[10][6],pp[9][7],pp[8][8],s_0_16_7,c_0_16_7);
    wire s_0_16_8, c_0_16_8;
    csa u_csa_0_16_8(pp[7][9],pp[6][10],pp[5][11],s_0_16_8,c_0_16_8);
    wire s_0_16_9, c_0_16_9;
    csa u_csa_0_16_9(pp[4][12],pp[3][13],pp[2][14],s_0_16_9,c_0_16_9);
    wire s_0_17_5, c_0_17_5;
    csa u_csa_0_17_5(pp[17][0],pp[16][1],pp[15][2],s_0_17_5,c_0_17_5);
    wire s_0_17_6, c_0_17_6;
    csa u_csa_0_17_6(pp[14][3],pp[13][4],pp[12][5],s_0_17_6,c_0_17_6);
    wire s_0_17_7, c_0_17_7;
    csa u_csa_0_17_7(pp[11][6],pp[10][7],pp[9][8],s_0_17_7,c_0_17_7);
    wire s_0_17_8, c_0_17_8;
    csa u_csa_0_17_8(pp[8][9],pp[7][10],pp[6][11],s_0_17_8,c_0_17_8);
    wire s_0_17_9, c_0_17_9;
    csa u_csa_0_17_9(pp[5][12],pp[4][13],pp[3][14],s_0_17_9,c_0_17_9);
    wire s_0_17_10, c_0_17_10;
    csa u_csa_0_17_10(pp[2][15],pp[1][16],pp[0][17],s_0_17_10,c_0_17_10);
    wire s_0_18_6, c_0_18_6;
    csa u_csa_0_18_6(pp[18][0],pp[17][1],pp[16][2],s_0_18_6,c_0_18_6);
    wire s_0_18_7, c_0_18_7;
    csa u_csa_0_18_7(pp[15][3],pp[14][4],pp[13][5],s_0_18_7,c_0_18_7);
    wire s_0_18_8, c_0_18_8;
    csa u_csa_0_18_8(pp[12][6],pp[11][7],pp[10][8],s_0_18_8,c_0_18_8);
    wire s_0_18_9, c_0_18_9;
    csa u_csa_0_18_9(pp[9][9],pp[8][10],pp[7][11],s_0_18_9,c_0_18_9);
    wire s_0_18_10, c_0_18_10;
    csa u_csa_0_18_10(pp[6][12],pp[5][13],pp[4][14],s_0_18_10,c_0_18_10);
    wire s_0_18_11, c_0_18_11;
    csa u_csa_0_18_11(pp[3][15],pp[2][16],pp[1][17],s_0_18_11,c_0_18_11);
    wire s_0_19_6, c_0_19_6;
    csa u_csa_0_19_6(pp[19][0],pp[18][1],pp[17][2],s_0_19_6,c_0_19_6);
    wire s_0_19_7, c_0_19_7;
    csa u_csa_0_19_7(pp[16][3],pp[15][4],pp[14][5],s_0_19_7,c_0_19_7);
    wire s_0_19_8, c_0_19_8;
    csa u_csa_0_19_8(pp[13][6],pp[12][7],pp[11][8],s_0_19_8,c_0_19_8);
    wire s_0_19_9, c_0_19_9;
    csa u_csa_0_19_9(pp[10][9],pp[9][10],pp[8][11],s_0_19_9,c_0_19_9);
    wire s_0_19_10, c_0_19_10;
    csa u_csa_0_19_10(pp[7][12],pp[6][13],pp[5][14],s_0_19_10,c_0_19_10);
    wire s_0_19_11, c_0_19_11;
    csa u_csa_0_19_11(pp[4][15],pp[3][16],pp[2][17],s_0_19_11,c_0_19_11);
    wire s_0_20_6, c_0_20_6;
    csa u_csa_0_20_6(pp[20][0],pp[19][1],pp[18][2],s_0_20_6,c_0_20_6);
    wire s_0_20_7, c_0_20_7;
    csa u_csa_0_20_7(pp[17][3],pp[16][4],pp[15][5],s_0_20_7,c_0_20_7);
    wire s_0_20_8, c_0_20_8;
    csa u_csa_0_20_8(pp[14][6],pp[13][7],pp[12][8],s_0_20_8,c_0_20_8);
    wire s_0_20_9, c_0_20_9;
    csa u_csa_0_20_9(pp[11][9],pp[10][10],pp[9][11],s_0_20_9,c_0_20_9);
    wire s_0_20_10, c_0_20_10;
    csa u_csa_0_20_10(pp[8][12],pp[7][13],pp[6][14],s_0_20_10,c_0_20_10);
    wire s_0_20_11, c_0_20_11;
    csa u_csa_0_20_11(pp[5][15],pp[4][16],pp[3][17],s_0_20_11,c_0_20_11);
    wire s_0_20_12, c_0_20_12;
    csa u_csa_0_20_12(pp[2][18],pp[1][19],pp[0][20],s_0_20_12,c_0_20_12);
    wire s_0_21_7, c_0_21_7;
    csa u_csa_0_21_7(pp[21][0],pp[20][1],pp[19][2],s_0_21_7,c_0_21_7);
    wire s_0_21_8, c_0_21_8;
    csa u_csa_0_21_8(pp[18][3],pp[17][4],pp[16][5],s_0_21_8,c_0_21_8);
    wire s_0_21_9, c_0_21_9;
    csa u_csa_0_21_9(pp[15][6],pp[14][7],pp[13][8],s_0_21_9,c_0_21_9);
    wire s_0_21_10, c_0_21_10;
    csa u_csa_0_21_10(pp[12][9],pp[11][10],pp[10][11],s_0_21_10,c_0_21_10);
    wire s_0_21_11, c_0_21_11;
    csa u_csa_0_21_11(pp[9][12],pp[8][13],pp[7][14],s_0_21_11,c_0_21_11);
    wire s_0_21_12, c_0_21_12;
    csa u_csa_0_21_12(pp[6][15],pp[5][16],pp[4][17],s_0_21_12,c_0_21_12);
    wire s_0_21_13, c_0_21_13;
    csa u_csa_0_21_13(pp[3][18],pp[2][19],pp[1][20],s_0_21_13,c_0_21_13);
    wire s_0_22_7, c_0_22_7;
    csa u_csa_0_22_7(pp[22][0],pp[21][1],pp[20][2],s_0_22_7,c_0_22_7);
    wire s_0_22_8, c_0_22_8;
    csa u_csa_0_22_8(pp[19][3],pp[18][4],pp[17][5],s_0_22_8,c_0_22_8);
    wire s_0_22_9, c_0_22_9;
    csa u_csa_0_22_9(pp[16][6],pp[15][7],pp[14][8],s_0_22_9,c_0_22_9);
    wire s_0_22_10, c_0_22_10;
    csa u_csa_0_22_10(pp[13][9],pp[12][10],pp[11][11],s_0_22_10,c_0_22_10);
    wire s_0_22_11, c_0_22_11;
    csa u_csa_0_22_11(pp[10][12],pp[9][13],pp[8][14],s_0_22_11,c_0_22_11);
    wire s_0_22_12, c_0_22_12;
    csa u_csa_0_22_12(pp[7][15],pp[6][16],pp[5][17],s_0_22_12,c_0_22_12);
    wire s_0_22_13, c_0_22_13;
    csa u_csa_0_22_13(pp[4][18],pp[3][19],pp[2][20],s_0_22_13,c_0_22_13);
    wire s_0_23_7, c_0_23_7;
    csa u_csa_0_23_7(pp[23][0],pp[22][1],pp[21][2],s_0_23_7,c_0_23_7);
    wire s_0_23_8, c_0_23_8;
    csa u_csa_0_23_8(pp[20][3],pp[19][4],pp[18][5],s_0_23_8,c_0_23_8);
    wire s_0_23_9, c_0_23_9;
    csa u_csa_0_23_9(pp[17][6],pp[16][7],pp[15][8],s_0_23_9,c_0_23_9);
    wire s_0_23_10, c_0_23_10;
    csa u_csa_0_23_10(pp[14][9],pp[13][10],pp[12][11],s_0_23_10,c_0_23_10);
    wire s_0_23_11, c_0_23_11;
    csa u_csa_0_23_11(pp[11][12],pp[10][13],pp[9][14],s_0_23_11,c_0_23_11);
    wire s_0_23_12, c_0_23_12;
    csa u_csa_0_23_12(pp[8][15],pp[7][16],pp[6][17],s_0_23_12,c_0_23_12);
    wire s_0_23_13, c_0_23_13;
    csa u_csa_0_23_13(pp[5][18],pp[4][19],pp[3][20],s_0_23_13,c_0_23_13);
    wire s_0_23_14, c_0_23_14;
    csa u_csa_0_23_14(pp[2][21],pp[1][22],pp[0][23],s_0_23_14,c_0_23_14);
    wire s_0_24_8, c_0_24_8;
    csa u_csa_0_24_8(pp[24][0],pp[23][1],pp[22][2],s_0_24_8,c_0_24_8);
    wire s_0_24_9, c_0_24_9;
    csa u_csa_0_24_9(pp[21][3],pp[20][4],pp[19][5],s_0_24_9,c_0_24_9);
    wire s_0_24_10, c_0_24_10;
    csa u_csa_0_24_10(pp[18][6],pp[17][7],pp[16][8],s_0_24_10,c_0_24_10);
    wire s_0_24_11, c_0_24_11;
    csa u_csa_0_24_11(pp[15][9],pp[14][10],pp[13][11],s_0_24_11,c_0_24_11);
    wire s_0_24_12, c_0_24_12;
    csa u_csa_0_24_12(pp[12][12],pp[11][13],pp[10][14],s_0_24_12,c_0_24_12);
    wire s_0_24_13, c_0_24_13;
    csa u_csa_0_24_13(pp[9][15],pp[8][16],pp[7][17],s_0_24_13,c_0_24_13);
    wire s_0_24_14, c_0_24_14;
    csa u_csa_0_24_14(pp[6][18],pp[5][19],pp[4][20],s_0_24_14,c_0_24_14);
    wire s_0_24_15, c_0_24_15;
    csa u_csa_0_24_15(pp[3][21],pp[2][22],pp[1][23],s_0_24_15,c_0_24_15);
    wire s_0_25_8, c_0_25_8;
    csa u_csa_0_25_8(pp[25][0],pp[24][1],pp[23][2],s_0_25_8,c_0_25_8);
    wire s_0_25_9, c_0_25_9;
    csa u_csa_0_25_9(pp[22][3],pp[21][4],pp[20][5],s_0_25_9,c_0_25_9);
    wire s_0_25_10, c_0_25_10;
    csa u_csa_0_25_10(pp[19][6],pp[18][7],pp[17][8],s_0_25_10,c_0_25_10);
    wire s_0_25_11, c_0_25_11;
    csa u_csa_0_25_11(pp[16][9],pp[15][10],pp[14][11],s_0_25_11,c_0_25_11);
    wire s_0_25_12, c_0_25_12;
    csa u_csa_0_25_12(pp[13][12],pp[12][13],pp[11][14],s_0_25_12,c_0_25_12);
    wire s_0_25_13, c_0_25_13;
    csa u_csa_0_25_13(pp[10][15],pp[9][16],pp[8][17],s_0_25_13,c_0_25_13);
    wire s_0_25_14, c_0_25_14;
    csa u_csa_0_25_14(pp[7][18],pp[6][19],pp[5][20],s_0_25_14,c_0_25_14);
    wire s_0_25_15, c_0_25_15;
    csa u_csa_0_25_15(pp[4][21],pp[3][22],pp[2][23],s_0_25_15,c_0_25_15);
    wire s_0_26_8, c_0_26_8;
    csa u_csa_0_26_8(pp[25][1],pp[24][2],pp[23][3],s_0_26_8,c_0_26_8);
    wire s_0_26_9, c_0_26_9;
    csa u_csa_0_26_9(pp[22][4],pp[21][5],pp[20][6],s_0_26_9,c_0_26_9);
    wire s_0_26_10, c_0_26_10;
    csa u_csa_0_26_10(pp[19][7],pp[18][8],pp[17][9],s_0_26_10,c_0_26_10);
    wire s_0_26_11, c_0_26_11;
    csa u_csa_0_26_11(pp[16][10],pp[15][11],pp[14][12],s_0_26_11,c_0_26_11);
    wire s_0_26_12, c_0_26_12;
    csa u_csa_0_26_12(pp[13][13],pp[12][14],pp[11][15],s_0_26_12,c_0_26_12);
    wire s_0_26_13, c_0_26_13;
    csa u_csa_0_26_13(pp[10][16],pp[9][17],pp[8][18],s_0_26_13,c_0_26_13);
    wire s_0_26_14, c_0_26_14;
    csa u_csa_0_26_14(pp[7][19],pp[6][20],pp[5][21],s_0_26_14,c_0_26_14);
    wire s_0_26_15, c_0_26_15;
    csa u_csa_0_26_15(pp[4][22],pp[3][23],pp[2][24],s_0_26_15,c_0_26_15);
    wire s_0_27_8, c_0_27_8;
    csa u_csa_0_27_8(pp[25][2],pp[24][3],pp[23][4],s_0_27_8,c_0_27_8);
    wire s_0_27_9, c_0_27_9;
    csa u_csa_0_27_9(pp[22][5],pp[21][6],pp[20][7],s_0_27_9,c_0_27_9);
    wire s_0_27_10, c_0_27_10;
    csa u_csa_0_27_10(pp[19][8],pp[18][9],pp[17][10],s_0_27_10,c_0_27_10);
    wire s_0_27_11, c_0_27_11;
    csa u_csa_0_27_11(pp[16][11],pp[15][12],pp[14][13],s_0_27_11,c_0_27_11);
    wire s_0_27_12, c_0_27_12;
    csa u_csa_0_27_12(pp[13][14],pp[12][15],pp[11][16],s_0_27_12,c_0_27_12);
    wire s_0_27_13, c_0_27_13;
    csa u_csa_0_27_13(pp[10][17],pp[9][18],pp[8][19],s_0_27_13,c_0_27_13);
    wire s_0_27_14, c_0_27_14;
    csa u_csa_0_27_14(pp[7][20],pp[6][21],pp[5][22],s_0_27_14,c_0_27_14);
    wire s_0_27_15, c_0_27_15;
    csa u_csa_0_27_15(pp[4][23],pp[3][24],pp[2][25],s_0_27_15,c_0_27_15);
    wire s_0_28_8, c_0_28_8;
    csa u_csa_0_28_8(pp[25][3],pp[24][4],pp[23][5],s_0_28_8,c_0_28_8);
    wire s_0_28_9, c_0_28_9;
    csa u_csa_0_28_9(pp[22][6],pp[21][7],pp[20][8],s_0_28_9,c_0_28_9);
    wire s_0_28_10, c_0_28_10;
    csa u_csa_0_28_10(pp[19][9],pp[18][10],pp[17][11],s_0_28_10,c_0_28_10);
    wire s_0_28_11, c_0_28_11;
    csa u_csa_0_28_11(pp[16][12],pp[15][13],pp[14][14],s_0_28_11,c_0_28_11);
    wire s_0_28_12, c_0_28_12;
    csa u_csa_0_28_12(pp[13][15],pp[12][16],pp[11][17],s_0_28_12,c_0_28_12);
    wire s_0_28_13, c_0_28_13;
    csa u_csa_0_28_13(pp[10][18],pp[9][19],pp[8][20],s_0_28_13,c_0_28_13);
    wire s_0_28_14, c_0_28_14;
    csa u_csa_0_28_14(pp[7][21],pp[6][22],pp[5][23],s_0_28_14,c_0_28_14);
    wire s_0_29_7, c_0_29_7;
    csa u_csa_0_29_7(pp[25][4],pp[24][5],pp[23][6],s_0_29_7,c_0_29_7);
    wire s_0_29_8, c_0_29_8;
    csa u_csa_0_29_8(pp[22][7],pp[21][8],pp[20][9],s_0_29_8,c_0_29_8);
    wire s_0_29_9, c_0_29_9;
    csa u_csa_0_29_9(pp[19][10],pp[18][11],pp[17][12],s_0_29_9,c_0_29_9);
    wire s_0_29_10, c_0_29_10;
    csa u_csa_0_29_10(pp[16][13],pp[15][14],pp[14][15],s_0_29_10,c_0_29_10);
    wire s_0_29_11, c_0_29_11;
    csa u_csa_0_29_11(pp[13][16],pp[12][17],pp[11][18],s_0_29_11,c_0_29_11);
    wire s_0_29_12, c_0_29_12;
    csa u_csa_0_29_12(pp[10][19],pp[9][20],pp[8][21],s_0_29_12,c_0_29_12);
    wire s_0_29_13, c_0_29_13;
    csa u_csa_0_29_13(pp[7][22],pp[6][23],pp[5][24],s_0_29_13,c_0_29_13);
    wire s_0_30_7, c_0_30_7;
    csa u_csa_0_30_7(pp[25][5],pp[24][6],pp[23][7],s_0_30_7,c_0_30_7);
    wire s_0_30_8, c_0_30_8;
    csa u_csa_0_30_8(pp[22][8],pp[21][9],pp[20][10],s_0_30_8,c_0_30_8);
    wire s_0_30_9, c_0_30_9;
    csa u_csa_0_30_9(pp[19][11],pp[18][12],pp[17][13],s_0_30_9,c_0_30_9);
    wire s_0_30_10, c_0_30_10;
    csa u_csa_0_30_10(pp[16][14],pp[15][15],pp[14][16],s_0_30_10,c_0_30_10);
    wire s_0_30_11, c_0_30_11;
    csa u_csa_0_30_11(pp[13][17],pp[12][18],pp[11][19],s_0_30_11,c_0_30_11);
    wire s_0_30_12, c_0_30_12;
    csa u_csa_0_30_12(pp[10][20],pp[9][21],pp[8][22],s_0_30_12,c_0_30_12);
    wire s_0_30_13, c_0_30_13;
    csa u_csa_0_30_13(pp[7][23],pp[6][24],pp[5][25],s_0_30_13,c_0_30_13);
    wire s_0_31_7, c_0_31_7;
    csa u_csa_0_31_7(pp[25][6],pp[24][7],pp[23][8],s_0_31_7,c_0_31_7);
    wire s_0_31_8, c_0_31_8;
    csa u_csa_0_31_8(pp[22][9],pp[21][10],pp[20][11],s_0_31_8,c_0_31_8);
    wire s_0_31_9, c_0_31_9;
    csa u_csa_0_31_9(pp[19][12],pp[18][13],pp[17][14],s_0_31_9,c_0_31_9);
    wire s_0_31_10, c_0_31_10;
    csa u_csa_0_31_10(pp[16][15],pp[15][16],pp[14][17],s_0_31_10,c_0_31_10);
    wire s_0_31_11, c_0_31_11;
    csa u_csa_0_31_11(pp[13][18],pp[12][19],pp[11][20],s_0_31_11,c_0_31_11);
    wire s_0_31_12, c_0_31_12;
    csa u_csa_0_31_12(pp[10][21],pp[9][22],pp[8][23],s_0_31_12,c_0_31_12);
    wire s_0_32_6, c_0_32_6;
    csa u_csa_0_32_6(pp[25][7],pp[24][8],pp[23][9],s_0_32_6,c_0_32_6);
    wire s_0_32_7, c_0_32_7;
    csa u_csa_0_32_7(pp[22][10],pp[21][11],pp[20][12],s_0_32_7,c_0_32_7);
    wire s_0_32_8, c_0_32_8;
    csa u_csa_0_32_8(pp[19][13],pp[18][14],pp[17][15],s_0_32_8,c_0_32_8);
    wire s_0_32_9, c_0_32_9;
    csa u_csa_0_32_9(pp[16][16],pp[15][17],pp[14][18],s_0_32_9,c_0_32_9);
    wire s_0_32_10, c_0_32_10;
    csa u_csa_0_32_10(pp[13][19],pp[12][20],pp[11][21],s_0_32_10,c_0_32_10);
    wire s_0_32_11, c_0_32_11;
    csa u_csa_0_32_11(pp[10][22],pp[9][23],pp[8][24],s_0_32_11,c_0_32_11);
    wire s_0_33_6, c_0_33_6;
    csa u_csa_0_33_6(pp[25][8],pp[24][9],pp[23][10],s_0_33_6,c_0_33_6);
    wire s_0_33_7, c_0_33_7;
    csa u_csa_0_33_7(pp[22][11],pp[21][12],pp[20][13],s_0_33_7,c_0_33_7);
    wire s_0_33_8, c_0_33_8;
    csa u_csa_0_33_8(pp[19][14],pp[18][15],pp[17][16],s_0_33_8,c_0_33_8);
    wire s_0_33_9, c_0_33_9;
    csa u_csa_0_33_9(pp[16][17],pp[15][18],pp[14][19],s_0_33_9,c_0_33_9);
    wire s_0_33_10, c_0_33_10;
    csa u_csa_0_33_10(pp[13][20],pp[12][21],pp[11][22],s_0_33_10,c_0_33_10);
    wire s_0_33_11, c_0_33_11;
    csa u_csa_0_33_11(pp[10][23],pp[9][24],pp[8][25],s_0_33_11,c_0_33_11);
    wire s_0_34_6, c_0_34_6;
    csa u_csa_0_34_6(pp[25][9],pp[24][10],pp[23][11],s_0_34_6,c_0_34_6);
    wire s_0_34_7, c_0_34_7;
    csa u_csa_0_34_7(pp[22][12],pp[21][13],pp[20][14],s_0_34_7,c_0_34_7);
    wire s_0_34_8, c_0_34_8;
    csa u_csa_0_34_8(pp[19][15],pp[18][16],pp[17][17],s_0_34_8,c_0_34_8);
    wire s_0_34_9, c_0_34_9;
    csa u_csa_0_34_9(pp[16][18],pp[15][19],pp[14][20],s_0_34_9,c_0_34_9);
    wire s_0_34_10, c_0_34_10;
    csa u_csa_0_34_10(pp[13][21],pp[12][22],pp[11][23],s_0_34_10,c_0_34_10);
    wire s_0_35_5, c_0_35_5;
    csa u_csa_0_35_5(pp[25][10],pp[24][11],pp[23][12],s_0_35_5,c_0_35_5);
    wire s_0_35_6, c_0_35_6;
    csa u_csa_0_35_6(pp[22][13],pp[21][14],pp[20][15],s_0_35_6,c_0_35_6);
    wire s_0_35_7, c_0_35_7;
    csa u_csa_0_35_7(pp[19][16],pp[18][17],pp[17][18],s_0_35_7,c_0_35_7);
    wire s_0_35_8, c_0_35_8;
    csa u_csa_0_35_8(pp[16][19],pp[15][20],pp[14][21],s_0_35_8,c_0_35_8);
    wire s_0_35_9, c_0_35_9;
    csa u_csa_0_35_9(pp[13][22],pp[12][23],pp[11][24],s_0_35_9,c_0_35_9);
    wire s_0_36_5, c_0_36_5;
    csa u_csa_0_36_5(pp[25][11],pp[24][12],pp[23][13],s_0_36_5,c_0_36_5);
    wire s_0_36_6, c_0_36_6;
    csa u_csa_0_36_6(pp[22][14],pp[21][15],pp[20][16],s_0_36_6,c_0_36_6);
    wire s_0_36_7, c_0_36_7;
    csa u_csa_0_36_7(pp[19][17],pp[18][18],pp[17][19],s_0_36_7,c_0_36_7);
    wire s_0_36_8, c_0_36_8;
    csa u_csa_0_36_8(pp[16][20],pp[15][21],pp[14][22],s_0_36_8,c_0_36_8);
    wire s_0_36_9, c_0_36_9;
    csa u_csa_0_36_9(pp[13][23],pp[12][24],pp[11][25],s_0_36_9,c_0_36_9);
    wire s_0_37_5, c_0_37_5;
    csa u_csa_0_37_5(pp[25][12],pp[24][13],pp[23][14],s_0_37_5,c_0_37_5);
    wire s_0_37_6, c_0_37_6;
    csa u_csa_0_37_6(pp[22][15],pp[21][16],pp[20][17],s_0_37_6,c_0_37_6);
    wire s_0_37_7, c_0_37_7;
    csa u_csa_0_37_7(pp[19][18],pp[18][19],pp[17][20],s_0_37_7,c_0_37_7);
    wire s_0_37_8, c_0_37_8;
    csa u_csa_0_37_8(pp[16][21],pp[15][22],pp[14][23],s_0_37_8,c_0_37_8);
    wire s_0_38_4, c_0_38_4;
    csa u_csa_0_38_4(pp[25][13],pp[24][14],pp[23][15],s_0_38_4,c_0_38_4);
    wire s_0_38_5, c_0_38_5;
    csa u_csa_0_38_5(pp[22][16],pp[21][17],pp[20][18],s_0_38_5,c_0_38_5);
    wire s_0_38_6, c_0_38_6;
    csa u_csa_0_38_6(pp[19][19],pp[18][20],pp[17][21],s_0_38_6,c_0_38_6);
    wire s_0_38_7, c_0_38_7;
    csa u_csa_0_38_7(pp[16][22],pp[15][23],pp[14][24],s_0_38_7,c_0_38_7);
    wire s_0_39_4, c_0_39_4;
    csa u_csa_0_39_4(pp[25][14],pp[24][15],pp[23][16],s_0_39_4,c_0_39_4);
    wire s_0_39_5, c_0_39_5;
    csa u_csa_0_39_5(pp[22][17],pp[21][18],pp[20][19],s_0_39_5,c_0_39_5);
    wire s_0_39_6, c_0_39_6;
    csa u_csa_0_39_6(pp[19][20],pp[18][21],pp[17][22],s_0_39_6,c_0_39_6);
    wire s_0_39_7, c_0_39_7;
    csa u_csa_0_39_7(pp[16][23],pp[15][24],pp[14][25],s_0_39_7,c_0_39_7);
    wire s_0_40_4, c_0_40_4;
    csa u_csa_0_40_4(pp[25][15],pp[24][16],pp[23][17],s_0_40_4,c_0_40_4);
    wire s_0_40_5, c_0_40_5;
    csa u_csa_0_40_5(pp[22][18],pp[21][19],pp[20][20],s_0_40_5,c_0_40_5);
    wire s_0_40_6, c_0_40_6;
    csa u_csa_0_40_6(pp[19][21],pp[18][22],pp[17][23],s_0_40_6,c_0_40_6);
    wire s_0_41_3, c_0_41_3;
    csa u_csa_0_41_3(pp[25][16],pp[24][17],pp[23][18],s_0_41_3,c_0_41_3);
    wire s_0_41_4, c_0_41_4;
    csa u_csa_0_41_4(pp[22][19],pp[21][20],pp[20][21],s_0_41_4,c_0_41_4);
    wire s_0_41_5, c_0_41_5;
    csa u_csa_0_41_5(pp[19][22],pp[18][23],pp[17][24],s_0_41_5,c_0_41_5);
    wire s_0_42_3, c_0_42_3;
    csa u_csa_0_42_3(pp[25][17],pp[24][18],pp[23][19],s_0_42_3,c_0_42_3);
    wire s_0_42_4, c_0_42_4;
    csa u_csa_0_42_4(pp[22][20],pp[21][21],pp[20][22],s_0_42_4,c_0_42_4);
    wire s_0_42_5, c_0_42_5;
    csa u_csa_0_42_5(pp[19][23],pp[18][24],pp[17][25],s_0_42_5,c_0_42_5);
    wire s_0_43_3, c_0_43_3;
    csa u_csa_0_43_3(pp[25][18],pp[24][19],pp[23][20],s_0_43_3,c_0_43_3);
    wire s_0_43_4, c_0_43_4;
    csa u_csa_0_43_4(pp[22][21],pp[21][22],pp[20][23],s_0_43_4,c_0_43_4);
    wire s_0_44_2, c_0_44_2;
    csa u_csa_0_44_2(pp[25][19],pp[24][20],pp[23][21],s_0_44_2,c_0_44_2);
    wire s_0_44_3, c_0_44_3;
    csa u_csa_0_44_3(pp[22][22],pp[21][23],pp[20][24],s_0_44_3,c_0_44_3);
    wire s_0_45_2, c_0_45_2;
    csa u_csa_0_45_2(pp[25][20],pp[24][21],pp[23][22],s_0_45_2,c_0_45_2);
    wire s_0_45_3, c_0_45_3;
    csa u_csa_0_45_3(pp[22][23],pp[21][24],pp[20][25],s_0_45_3,c_0_45_3);
    wire s_0_46_2, c_0_46_2;
    csa u_csa_0_46_2(pp[25][21],pp[24][22],pp[23][23],s_0_46_2,c_0_46_2);
    wire s_0_47_1, c_0_47_1;
    csa u_csa_0_47_1(pp[25][22],pp[24][23],pp[23][24],s_0_47_1,c_0_47_1);
    wire s_0_48_1, c_0_48_1;
    csa u_csa_0_48_1(pp[25][23],pp[24][24],pp[23][25],s_0_48_1,c_0_48_1);
    wire s_1_3_0, c_1_3_0;
    csa u_csa_1_3_0(pp[0][3],s_0_3_1,c_0_2_0,s_1_3_0,c_1_3_0);
    wire s_1_4_1, c_1_4_1;
    csa u_csa_1_4_1(pp[0][4],pp[1][3],s_0_4_1,s_1_4_1,c_1_4_1);
    wire s_1_5_1, c_1_5_1;
    csa u_csa_1_5_1(s_0_5_2,s_0_5_1,c_0_4_1,s_1_5_1,c_1_5_1);
    wire s_1_6_1, c_1_6_1;
    csa u_csa_1_6_1(pp[0][6],s_0_6_3,s_0_6_2,s_1_6_1,c_1_6_1);
    wire s_1_7_1, c_1_7_1;
    csa u_csa_1_7_1(pp[0][7],pp[1][6],s_0_7_3,s_1_7_1,c_1_7_1);
    wire s_1_7_2, c_1_7_2;
    csa u_csa_1_7_2(s_0_7_2,c_0_6_3,c_0_6_2,s_1_7_2,c_1_7_2);
    wire s_1_8_2, c_1_8_2;
    csa u_csa_1_8_2(s_0_8_4,s_0_8_3,s_0_8_2,s_1_8_2,c_1_8_2);
    wire s_1_9_1, c_1_9_1;
    csa u_csa_1_9_1(pp[0][9],s_0_9_5,s_0_9_4,s_1_9_1,c_1_9_1);
    wire s_1_9_2, c_1_9_2;
    csa u_csa_1_9_2(s_0_9_3,c_0_8_4,c_0_8_3,s_1_9_2,c_1_9_2);
    wire s_1_10_2, c_1_10_2;
    csa u_csa_1_10_2(pp[0][10],pp[1][9],s_0_10_5,s_1_10_2,c_1_10_2);
    wire s_1_10_3, c_1_10_3;
    csa u_csa_1_10_3(s_0_10_4,s_0_10_3,c_0_9_5,s_1_10_3,c_1_10_3);
    wire s_1_11_2, c_1_11_2;
    csa u_csa_1_11_2(s_0_11_6,s_0_11_5,s_0_11_4,s_1_11_2,c_1_11_2);
    wire s_1_11_3, c_1_11_3;
    csa u_csa_1_11_3(s_0_11_3,c_0_10_5,c_0_10_4,s_1_11_3,c_1_11_3);
    wire s_1_12_2, c_1_12_2;
    csa u_csa_1_12_2(pp[0][12],s_0_12_7,s_0_12_6,s_1_12_2,c_1_12_2);
    wire s_1_12_3, c_1_12_3;
    csa u_csa_1_12_3(s_0_12_5,s_0_12_4,c_0_11_6,s_1_12_3,c_1_12_3);
    wire s_1_12_4, c_1_12_4;
    csa u_csa_1_12_4(c_0_11_5,c_0_11_4,c_0_11_3,s_1_12_4,c_1_12_4);
    wire s_1_13_3, c_1_13_3;
    csa u_csa_1_13_3(pp[0][13],pp[1][12],s_0_13_7,s_1_13_3,c_1_13_3);
    wire s_1_13_4, c_1_13_4;
    csa u_csa_1_13_4(s_0_13_6,s_0_13_5,s_0_13_4,s_1_13_4,c_1_13_4);
    wire s_1_13_5, c_1_13_5;
    csa u_csa_1_13_5(c_0_12_7,c_0_12_6,c_0_12_5,s_1_13_5,c_1_13_5);
    wire s_1_14_3, c_1_14_3;
    csa u_csa_1_14_3(s_0_14_8,s_0_14_7,s_0_14_6,s_1_14_3,c_1_14_3);
    wire s_1_14_4, c_1_14_4;
    csa u_csa_1_14_4(s_0_14_5,s_0_14_4,c_0_13_7,s_1_14_4,c_1_14_4);
    wire s_1_14_5, c_1_14_5;
    csa u_csa_1_14_5(c_0_13_6,c_0_13_5,c_0_13_4,s_1_14_5,c_1_14_5);
    wire s_1_15_3, c_1_15_3;
    csa u_csa_1_15_3(pp[0][15],s_0_15_9,s_0_15_8,s_1_15_3,c_1_15_3);
    wire s_1_15_4, c_1_15_4;
    csa u_csa_1_15_4(s_0_15_7,s_0_15_6,s_0_15_5,s_1_15_4,c_1_15_4);
    wire s_1_15_5, c_1_15_5;
    csa u_csa_1_15_5(c_0_14_8,c_0_14_7,c_0_14_6,s_1_15_5,c_1_15_5);
    wire s_1_16_3, c_1_16_3;
    csa u_csa_1_16_3(pp[0][16],pp[1][15],s_0_16_9,s_1_16_3,c_1_16_3);
    wire s_1_16_4, c_1_16_4;
    csa u_csa_1_16_4(s_0_16_8,s_0_16_7,s_0_16_6,s_1_16_4,c_1_16_4);
    wire s_1_16_5, c_1_16_5;
    csa u_csa_1_16_5(s_0_16_5,c_0_15_9,c_0_15_8,s_1_16_5,c_1_16_5);
    wire s_1_16_6, c_1_16_6;
    csa u_csa_1_16_6(c_0_15_7,c_0_15_6,c_0_15_5,s_1_16_6,c_1_16_6);
    wire s_1_17_4, c_1_17_4;
    csa u_csa_1_17_4(s_0_17_10,s_0_17_9,s_0_17_8,s_1_17_4,c_1_17_4);
    wire s_1_17_5, c_1_17_5;
    csa u_csa_1_17_5(s_0_17_7,s_0_17_6,s_0_17_5,s_1_17_5,c_1_17_5);
    wire s_1_17_6, c_1_17_6;
    csa u_csa_1_17_6(c_0_16_9,c_0_16_8,c_0_16_7,s_1_17_6,c_1_17_6);
    wire s_1_18_3, c_1_18_3;
    csa u_csa_1_18_3(pp[0][18],s_0_18_11,s_0_18_10,s_1_18_3,c_1_18_3);
    wire s_1_18_4, c_1_18_4;
    csa u_csa_1_18_4(s_0_18_9,s_0_18_8,s_0_18_7,s_1_18_4,c_1_18_4);
    wire s_1_18_5, c_1_18_5;
    csa u_csa_1_18_5(s_0_18_6,c_0_17_10,c_0_17_9,s_1_18_5,c_1_18_5);
    wire s_1_18_6, c_1_18_6;
    csa u_csa_1_18_6(c_0_17_8,c_0_17_7,c_0_17_6,s_1_18_6,c_1_18_6);
    wire s_1_19_4, c_1_19_4;
    csa u_csa_1_19_4(pp[0][19],pp[1][18],s_0_19_11,s_1_19_4,c_1_19_4);
    wire s_1_19_5, c_1_19_5;
    csa u_csa_1_19_5(s_0_19_10,s_0_19_9,s_0_19_8,s_1_19_5,c_1_19_5);
    wire s_1_19_6, c_1_19_6;
    csa u_csa_1_19_6(s_0_19_7,s_0_19_6,c_0_18_11,s_1_19_6,c_1_19_6);
    wire s_1_19_7, c_1_19_7;
    csa u_csa_1_19_7(c_0_18_10,c_0_18_9,c_0_18_8,s_1_19_7,c_1_19_7);
    wire s_1_20_4, c_1_20_4;
    csa u_csa_1_20_4(s_0_20_12,s_0_20_11,s_0_20_10,s_1_20_4,c_1_20_4);
    wire s_1_20_5, c_1_20_5;
    csa u_csa_1_20_5(s_0_20_9,s_0_20_8,s_0_20_7,s_1_20_5,c_1_20_5);
    wire s_1_20_6, c_1_20_6;
    csa u_csa_1_20_6(s_0_20_6,c_0_19_11,c_0_19_10,s_1_20_6,c_1_20_6);
    wire s_1_20_7, c_1_20_7;
    csa u_csa_1_20_7(c_0_19_9,c_0_19_8,c_0_19_7,s_1_20_7,c_1_20_7);
    wire s_1_21_4, c_1_21_4;
    csa u_csa_1_21_4(pp[0][21],s_0_21_13,s_0_21_12,s_1_21_4,c_1_21_4);
    wire s_1_21_5, c_1_21_5;
    csa u_csa_1_21_5(s_0_21_11,s_0_21_10,s_0_21_9,s_1_21_5,c_1_21_5);
    wire s_1_21_6, c_1_21_6;
    csa u_csa_1_21_6(s_0_21_8,s_0_21_7,c_0_20_12,s_1_21_6,c_1_21_6);
    wire s_1_21_7, c_1_21_7;
    csa u_csa_1_21_7(c_0_20_11,c_0_20_10,c_0_20_9,s_1_21_7,c_1_21_7);
    wire s_1_21_8, c_1_21_8;
    csa u_csa_1_21_8(c_0_20_8,c_0_20_7,c_0_20_6,s_1_21_8,c_1_21_8);
    wire s_1_22_5, c_1_22_5;
    csa u_csa_1_22_5(pp[0][22],pp[1][21],s_0_22_13,s_1_22_5,c_1_22_5);
    wire s_1_22_6, c_1_22_6;
    csa u_csa_1_22_6(s_0_22_12,s_0_22_11,s_0_22_10,s_1_22_6,c_1_22_6);
    wire s_1_22_7, c_1_22_7;
    csa u_csa_1_22_7(s_0_22_9,s_0_22_8,s_0_22_7,s_1_22_7,c_1_22_7);
    wire s_1_22_8, c_1_22_8;
    csa u_csa_1_22_8(c_0_21_13,c_0_21_12,c_0_21_11,s_1_22_8,c_1_22_8);
    wire s_1_22_9, c_1_22_9;
    csa u_csa_1_22_9(c_0_21_10,c_0_21_9,c_0_21_8,s_1_22_9,c_1_22_9);
    wire s_1_23_5, c_1_23_5;
    csa u_csa_1_23_5(s_0_23_14,s_0_23_13,s_0_23_12,s_1_23_5,c_1_23_5);
    wire s_1_23_6, c_1_23_6;
    csa u_csa_1_23_6(s_0_23_11,s_0_23_10,s_0_23_9,s_1_23_6,c_1_23_6);
    wire s_1_23_7, c_1_23_7;
    csa u_csa_1_23_7(s_0_23_8,s_0_23_7,c_0_22_13,s_1_23_7,c_1_23_7);
    wire s_1_23_8, c_1_23_8;
    csa u_csa_1_23_8(c_0_22_12,c_0_22_11,c_0_22_10,s_1_23_8,c_1_23_8);
    wire s_1_23_9, c_1_23_9;
    csa u_csa_1_23_9(c_0_22_9,c_0_22_8,c_0_22_7,s_1_23_9,c_1_23_9);
    wire s_1_24_5, c_1_24_5;
    csa u_csa_1_24_5(pp[0][24],s_0_24_15,s_0_24_14,s_1_24_5,c_1_24_5);
    wire s_1_24_6, c_1_24_6;
    csa u_csa_1_24_6(s_0_24_13,s_0_24_12,s_0_24_11,s_1_24_6,c_1_24_6);
    wire s_1_24_7, c_1_24_7;
    csa u_csa_1_24_7(s_0_24_10,s_0_24_9,s_0_24_8,s_1_24_7,c_1_24_7);
    wire s_1_24_8, c_1_24_8;
    csa u_csa_1_24_8(c_0_23_14,c_0_23_13,c_0_23_12,s_1_24_8,c_1_24_8);
    wire s_1_24_9, c_1_24_9;
    csa u_csa_1_24_9(c_0_23_11,c_0_23_10,c_0_23_9,s_1_24_9,c_1_24_9);
    wire s_1_25_5, c_1_25_5;
    csa u_csa_1_25_5(pp[0][25],pp[1][24],s_0_25_15,s_1_25_5,c_1_25_5);
    wire s_1_25_6, c_1_25_6;
    csa u_csa_1_25_6(s_0_25_14,s_0_25_13,s_0_25_12,s_1_25_6,c_1_25_6);
    wire s_1_25_7, c_1_25_7;
    csa u_csa_1_25_7(s_0_25_11,s_0_25_10,s_0_25_9,s_1_25_7,c_1_25_7);
    wire s_1_25_8, c_1_25_8;
    csa u_csa_1_25_8(s_0_25_8,c_0_24_15,c_0_24_14,s_1_25_8,c_1_25_8);
    wire s_1_25_9, c_1_25_9;
    csa u_csa_1_25_9(c_0_24_13,c_0_24_12,c_0_24_11,s_1_25_9,c_1_25_9);
    wire s_1_25_10, c_1_25_10;
    csa u_csa_1_25_10(c_0_24_10,c_0_24_9,c_0_24_8,s_1_25_10,c_1_25_10);
    wire s_1_26_6, c_1_26_6;
    csa u_csa_1_26_6(pp[1][25],s_0_26_15,s_0_26_14,s_1_26_6,c_1_26_6);
    wire s_1_26_7, c_1_26_7;
    csa u_csa_1_26_7(s_0_26_13,s_0_26_12,s_0_26_11,s_1_26_7,c_1_26_7);
    wire s_1_26_8, c_1_26_8;
    csa u_csa_1_26_8(s_0_26_10,s_0_26_9,s_0_26_8,s_1_26_8,c_1_26_8);
    wire s_1_26_9, c_1_26_9;
    csa u_csa_1_26_9(c_0_25_15,c_0_25_14,c_0_25_13,s_1_26_9,c_1_26_9);
    wire s_1_26_10, c_1_26_10;
    csa u_csa_1_26_10(c_0_25_12,c_0_25_11,c_0_25_10,s_1_26_10,c_1_26_10);
    wire s_1_27_5, c_1_27_5;
    csa u_csa_1_27_5(s_0_27_15,s_0_27_14,s_0_27_13,s_1_27_5,c_1_27_5);
    wire s_1_27_6, c_1_27_6;
    csa u_csa_1_27_6(s_0_27_12,s_0_27_11,s_0_27_10,s_1_27_6,c_1_27_6);
    wire s_1_27_7, c_1_27_7;
    csa u_csa_1_27_7(s_0_27_9,s_0_27_8,c_0_26_15,s_1_27_7,c_1_27_7);
    wire s_1_27_8, c_1_27_8;
    csa u_csa_1_27_8(c_0_26_14,c_0_26_13,c_0_26_12,s_1_27_8,c_1_27_8);
    wire s_1_27_9, c_1_27_9;
    csa u_csa_1_27_9(c_0_26_11,c_0_26_10,c_0_26_9,s_1_27_9,c_1_27_9);
    wire s_1_28_5, c_1_28_5;
    csa u_csa_1_28_5(pp[3][25],pp[4][24],s_0_28_14,s_1_28_5,c_1_28_5);
    wire s_1_28_6, c_1_28_6;
    csa u_csa_1_28_6(s_0_28_13,s_0_28_12,s_0_28_11,s_1_28_6,c_1_28_6);
    wire s_1_28_7, c_1_28_7;
    csa u_csa_1_28_7(s_0_28_10,s_0_28_9,s_0_28_8,s_1_28_7,c_1_28_7);
    wire s_1_28_8, c_1_28_8;
    csa u_csa_1_28_8(c_0_27_15,c_0_27_14,c_0_27_13,s_1_28_8,c_1_28_8);
    wire s_1_28_9, c_1_28_9;
    csa u_csa_1_28_9(c_0_27_12,c_0_27_11,c_0_27_10,s_1_28_9,c_1_28_9);
    wire s_1_29_5, c_1_29_5;
    csa u_csa_1_29_5(pp[4][25],s_0_29_13,s_0_29_12,s_1_29_5,c_1_29_5);
    wire s_1_29_6, c_1_29_6;
    csa u_csa_1_29_6(s_0_29_11,s_0_29_10,s_0_29_9,s_1_29_6,c_1_29_6);
    wire s_1_29_7, c_1_29_7;
    csa u_csa_1_29_7(s_0_29_8,s_0_29_7,c_0_28_14,s_1_29_7,c_1_29_7);
    wire s_1_29_8, c_1_29_8;
    csa u_csa_1_29_8(c_0_28_13,c_0_28_12,c_0_28_11,s_1_29_8,c_1_29_8);
    wire s_1_29_9, c_1_29_9;
    csa u_csa_1_29_9(c_0_28_10,c_0_28_9,c_0_28_8,s_1_29_9,c_1_29_9);
    wire s_1_30_5, c_1_30_5;
    csa u_csa_1_30_5(s_0_30_13,s_0_30_12,s_0_30_11,s_1_30_5,c_1_30_5);
    wire s_1_30_6, c_1_30_6;
    csa u_csa_1_30_6(s_0_30_10,s_0_30_9,s_0_30_8,s_1_30_6,c_1_30_6);
    wire s_1_30_7, c_1_30_7;
    csa u_csa_1_30_7(s_0_30_7,c_0_29_13,c_0_29_12,s_1_30_7,c_1_30_7);
    wire s_1_30_8, c_1_30_8;
    csa u_csa_1_30_8(c_0_29_11,c_0_29_10,c_0_29_9,s_1_30_8,c_1_30_8);
    wire s_1_31_4, c_1_31_4;
    csa u_csa_1_31_4(pp[6][25],pp[7][24],s_0_31_12,s_1_31_4,c_1_31_4);
    wire s_1_31_5, c_1_31_5;
    csa u_csa_1_31_5(s_0_31_11,s_0_31_10,s_0_31_9,s_1_31_5,c_1_31_5);
    wire s_1_31_6, c_1_31_6;
    csa u_csa_1_31_6(s_0_31_8,s_0_31_7,c_0_30_13,s_1_31_6,c_1_31_6);
    wire s_1_31_7, c_1_31_7;
    csa u_csa_1_31_7(c_0_30_12,c_0_30_11,c_0_30_10,s_1_31_7,c_1_31_7);
    wire s_1_31_8, c_1_31_8;
    csa u_csa_1_31_8(c_0_30_9,c_0_30_8,c_0_30_7,s_1_31_8,c_1_31_8);
    wire s_1_32_5, c_1_32_5;
    csa u_csa_1_32_5(pp[7][25],s_0_32_11,s_0_32_10,s_1_32_5,c_1_32_5);
    wire s_1_32_6, c_1_32_6;
    csa u_csa_1_32_6(s_0_32_9,s_0_32_8,s_0_32_7,s_1_32_6,c_1_32_6);
    wire s_1_32_7, c_1_32_7;
    csa u_csa_1_32_7(s_0_32_6,c_0_31_12,c_0_31_11,s_1_32_7,c_1_32_7);
    wire s_1_32_8, c_1_32_8;
    csa u_csa_1_32_8(c_0_31_10,c_0_31_9,c_0_31_8,s_1_32_8,c_1_32_8);
    wire s_1_33_4, c_1_33_4;
    csa u_csa_1_33_4(s_0_33_11,s_0_33_10,s_0_33_9,s_1_33_4,c_1_33_4);
    wire s_1_33_5, c_1_33_5;
    csa u_csa_1_33_5(s_0_33_8,s_0_33_7,s_0_33_6,s_1_33_5,c_1_33_5);
    wire s_1_33_6, c_1_33_6;
    csa u_csa_1_33_6(c_0_32_11,c_0_32_10,c_0_32_9,s_1_33_6,c_1_33_6);
    wire s_1_33_7, c_1_33_7;
    csa u_csa_1_33_7(c_0_32_8,c_0_32_7,c_0_32_6,s_1_33_7,c_1_33_7);
    wire s_1_34_4, c_1_34_4;
    csa u_csa_1_34_4(pp[9][25],pp[10][24],s_0_34_10,s_1_34_4,c_1_34_4);
    wire s_1_34_5, c_1_34_5;
    csa u_csa_1_34_5(s_0_34_9,s_0_34_8,s_0_34_7,s_1_34_5,c_1_34_5);
    wire s_1_34_6, c_1_34_6;
    csa u_csa_1_34_6(s_0_34_6,c_0_33_11,c_0_33_10,s_1_34_6,c_1_34_6);
    wire s_1_34_7, c_1_34_7;
    csa u_csa_1_34_7(c_0_33_9,c_0_33_8,c_0_33_7,s_1_34_7,c_1_34_7);
    wire s_1_35_4, c_1_35_4;
    csa u_csa_1_35_4(pp[10][25],s_0_35_9,s_0_35_8,s_1_35_4,c_1_35_4);
    wire s_1_35_5, c_1_35_5;
    csa u_csa_1_35_5(s_0_35_7,s_0_35_6,s_0_35_5,s_1_35_5,c_1_35_5);
    wire s_1_35_6, c_1_35_6;
    csa u_csa_1_35_6(c_0_34_10,c_0_34_9,c_0_34_8,s_1_35_6,c_1_35_6);
    wire s_1_36_3, c_1_36_3;
    csa u_csa_1_36_3(s_0_36_9,s_0_36_8,s_0_36_7,s_1_36_3,c_1_36_3);
    wire s_1_36_4, c_1_36_4;
    csa u_csa_1_36_4(s_0_36_6,s_0_36_5,c_0_35_9,s_1_36_4,c_1_36_4);
    wire s_1_36_5, c_1_36_5;
    csa u_csa_1_36_5(c_0_35_8,c_0_35_7,c_0_35_6,s_1_36_5,c_1_36_5);
    wire s_1_37_3, c_1_37_3;
    csa u_csa_1_37_3(pp[12][25],pp[13][24],s_0_37_8,s_1_37_3,c_1_37_3);
    wire s_1_37_4, c_1_37_4;
    csa u_csa_1_37_4(s_0_37_7,s_0_37_6,s_0_37_5,s_1_37_4,c_1_37_4);
    wire s_1_37_5, c_1_37_5;
    csa u_csa_1_37_5(c_0_36_9,c_0_36_8,c_0_36_7,s_1_37_5,c_1_37_5);
    wire s_1_38_3, c_1_38_3;
    csa u_csa_1_38_3(pp[13][25],s_0_38_7,s_0_38_6,s_1_38_3,c_1_38_3);
    wire s_1_38_4, c_1_38_4;
    csa u_csa_1_38_4(s_0_38_5,s_0_38_4,c_0_37_8,s_1_38_4,c_1_38_4);
    wire s_1_38_5, c_1_38_5;
    csa u_csa_1_38_5(c_0_37_7,c_0_37_6,c_0_37_5,s_1_38_5,c_1_38_5);
    wire s_1_39_3, c_1_39_3;
    csa u_csa_1_39_3(s_0_39_7,s_0_39_6,s_0_39_5,s_1_39_3,c_1_39_3);
    wire s_1_39_4, c_1_39_4;
    csa u_csa_1_39_4(s_0_39_4,c_0_38_7,c_0_38_6,s_1_39_4,c_1_39_4);
    wire s_1_40_2, c_1_40_2;
    csa u_csa_1_40_2(pp[15][25],pp[16][24],s_0_40_6,s_1_40_2,c_1_40_2);
    wire s_1_40_3, c_1_40_3;
    csa u_csa_1_40_3(s_0_40_5,s_0_40_4,c_0_39_7,s_1_40_3,c_1_40_3);
    wire s_1_40_4, c_1_40_4;
    csa u_csa_1_40_4(c_0_39_6,c_0_39_5,c_0_39_4,s_1_40_4,c_1_40_4);
    wire s_1_41_3, c_1_41_3;
    csa u_csa_1_41_3(pp[16][25],s_0_41_5,s_0_41_4,s_1_41_3,c_1_41_3);
    wire s_1_41_4, c_1_41_4;
    csa u_csa_1_41_4(s_0_41_3,c_0_40_6,c_0_40_5,s_1_41_4,c_1_41_4);
    wire s_1_42_2, c_1_42_2;
    csa u_csa_1_42_2(s_0_42_5,s_0_42_4,s_0_42_3,s_1_42_2,c_1_42_2);
    wire s_1_42_3, c_1_42_3;
    csa u_csa_1_42_3(c_0_41_5,c_0_41_4,c_0_41_3,s_1_42_3,c_1_42_3);
    wire s_1_43_2, c_1_43_2;
    csa u_csa_1_43_2(pp[18][25],pp[19][24],s_0_43_4,s_1_43_2,c_1_43_2);
    wire s_1_43_3, c_1_43_3;
    csa u_csa_1_43_3(s_0_43_3,c_0_42_5,c_0_42_4,s_1_43_3,c_1_43_3);
    wire s_1_44_2, c_1_44_2;
    csa u_csa_1_44_2(pp[19][25],s_0_44_3,s_0_44_2,s_1_44_2,c_1_44_2);
    wire s_1_45_1, c_1_45_1;
    csa u_csa_1_45_1(s_0_45_3,s_0_45_2,c_0_44_3,s_1_45_1,c_1_45_1);
    wire s_1_46_1, c_1_46_1;
    csa u_csa_1_46_1(pp[21][25],pp[22][24],s_0_46_2,s_1_46_1,c_1_46_1);
    wire s_1_47_1, c_1_47_1;
    csa u_csa_1_47_1(pp[22][25],s_0_47_1,c_0_46_2,s_1_47_1,c_1_47_1);
    wire s_1_49_0, c_1_49_0;
    csa u_csa_1_49_0(pp[24][25],pp[25][24],c_0_48_1,s_1_49_0,c_1_49_0);
    wire s_2_4_0, c_2_4_0;
    csa u_csa_2_4_0(c_0_3_1,s_1_4_1,c_1_3_0,s_2_4_0,c_2_4_0);
    wire s_2_6_0, c_2_6_0;
    csa u_csa_2_6_0(c_0_5_1,c_0_5_2,s_1_6_1,s_2_6_0,c_2_6_0);
    wire s_2_7_1, c_2_7_1;
    csa u_csa_2_7_1(s_1_7_2,s_1_7_1,c_1_6_1,s_2_7_1,c_2_7_1);
    wire s_2_8_1, c_2_8_1;
    csa u_csa_2_8_1(c_0_7_2,c_0_7_3,s_1_8_2,s_2_8_1,c_2_8_1);
    wire s_2_9_1, c_2_9_1;
    csa u_csa_2_9_1(c_0_8_2,s_1_9_2,s_1_9_1,s_2_9_1,c_2_9_1);
    wire s_2_10_1, c_2_10_1;
    csa u_csa_2_10_1(c_0_9_3,c_0_9_4,s_1_10_3,s_2_10_1,c_2_10_1);
    wire s_2_10_2, c_2_10_2;
    csa u_csa_2_10_2(s_1_10_2,c_1_9_2,c_1_9_1,s_2_10_2,c_2_10_2);
    wire s_2_11_2, c_2_11_2;
    csa u_csa_2_11_2(c_0_10_3,s_1_11_3,s_1_11_2,s_2_11_2,c_2_11_2);
    wire s_2_12_1, c_2_12_1;
    csa u_csa_2_12_1(s_1_12_4,s_1_12_3,s_1_12_2,s_2_12_1,c_2_12_1);
    wire s_2_13_1, c_2_13_1;
    csa u_csa_2_13_1(c_0_12_4,s_1_13_5,s_1_13_4,s_2_13_1,c_2_13_1);
    wire s_2_13_2, c_2_13_2;
    csa u_csa_2_13_2(s_1_13_3,c_1_12_4,c_1_12_3,s_2_13_2,c_2_13_2);
    wire s_2_14_2, c_2_14_2;
    csa u_csa_2_14_2(s_1_14_5,s_1_14_4,s_1_14_3,s_2_14_2,c_2_14_2);
    wire s_2_14_3, c_2_14_3;
    csa u_csa_2_14_3(c_1_13_5,c_1_13_4,c_1_13_3,s_2_14_3,c_2_14_3);
    wire s_2_15_2, c_2_15_2;
    csa u_csa_2_15_2(c_0_14_4,c_0_14_5,s_1_15_5,s_2_15_2,c_2_15_2);
    wire s_2_15_3, c_2_15_3;
    csa u_csa_2_15_3(s_1_15_4,s_1_15_3,c_1_14_5,s_2_15_3,c_2_15_3);
    wire s_2_16_2, c_2_16_2;
    csa u_csa_2_16_2(s_1_16_6,s_1_16_5,s_1_16_4,s_2_16_2,c_2_16_2);
    wire s_2_16_3, c_2_16_3;
    csa u_csa_2_16_3(s_1_16_3,c_1_15_5,c_1_15_4,s_2_16_3,c_2_16_3);
    wire s_2_17_2, c_2_17_2;
    csa u_csa_2_17_2(c_0_16_5,c_0_16_6,s_1_17_6,s_2_17_2,c_2_17_2);
    wire s_2_17_3, c_2_17_3;
    csa u_csa_2_17_3(s_1_17_5,s_1_17_4,c_1_16_6,s_2_17_3,c_2_17_3);
    wire s_2_17_4, c_2_17_4;
    csa u_csa_2_17_4(c_1_16_5,c_1_16_4,c_1_16_3,s_2_17_4,c_2_17_4);
    wire s_2_18_3, c_2_18_3;
    csa u_csa_2_18_3(c_0_17_5,s_1_18_6,s_1_18_5,s_2_18_3,c_2_18_3);
    wire s_2_18_4, c_2_18_4;
    csa u_csa_2_18_4(s_1_18_4,s_1_18_3,c_1_17_6,s_2_18_4,c_2_18_4);
    wire s_2_19_2, c_2_19_2;
    csa u_csa_2_19_2(c_0_18_6,c_0_18_7,s_1_19_7,s_2_19_2,c_2_19_2);
    wire s_2_19_3, c_2_19_3;
    csa u_csa_2_19_3(s_1_19_6,s_1_19_5,s_1_19_4,s_2_19_3,c_2_19_3);
    wire s_2_19_4, c_2_19_4;
    csa u_csa_2_19_4(c_1_18_6,c_1_18_5,c_1_18_4,s_2_19_4,c_2_19_4);
    wire s_2_20_3, c_2_20_3;
    csa u_csa_2_20_3(c_0_19_6,s_1_20_7,s_1_20_6,s_2_20_3,c_2_20_3);
    wire s_2_20_4, c_2_20_4;
    csa u_csa_2_20_4(s_1_20_5,s_1_20_4,c_1_19_7,s_2_20_4,c_2_20_4);
    wire s_2_20_5, c_2_20_5;
    csa u_csa_2_20_5(c_1_19_6,c_1_19_5,c_1_19_4,s_2_20_5,c_2_20_5);
    wire s_2_21_3, c_2_21_3;
    csa u_csa_2_21_3(s_1_21_8,s_1_21_7,s_1_21_6,s_2_21_3,c_2_21_3);
    wire s_2_21_4, c_2_21_4;
    csa u_csa_2_21_4(s_1_21_5,s_1_21_4,c_1_20_7,s_2_21_4,c_2_21_4);
    wire s_2_21_5, c_2_21_5;
    csa u_csa_2_21_5(c_1_20_6,c_1_20_5,c_1_20_4,s_2_21_5,c_2_21_5);
    wire s_2_22_3, c_2_22_3;
    csa u_csa_2_22_3(c_0_21_7,s_1_22_9,s_1_22_8,s_2_22_3,c_2_22_3);
    wire s_2_22_4, c_2_22_4;
    csa u_csa_2_22_4(s_1_22_7,s_1_22_6,s_1_22_5,s_2_22_4,c_2_22_4);
    wire s_2_22_5, c_2_22_5;
    csa u_csa_2_22_5(c_1_21_8,c_1_21_7,c_1_21_6,s_2_22_5,c_2_22_5);
    wire s_2_23_3, c_2_23_3;
    csa u_csa_2_23_3(s_1_23_9,s_1_23_8,s_1_23_7,s_2_23_3,c_2_23_3);
    wire s_2_23_4, c_2_23_4;
    csa u_csa_2_23_4(s_1_23_6,s_1_23_5,c_1_22_9,s_2_23_4,c_2_23_4);
    wire s_2_23_5, c_2_23_5;
    csa u_csa_2_23_5(c_1_22_8,c_1_22_7,c_1_22_6,s_2_23_5,c_2_23_5);
    wire s_2_24_3, c_2_24_3;
    csa u_csa_2_24_3(c_0_23_7,c_0_23_8,s_1_24_9,s_2_24_3,c_2_24_3);
    wire s_2_24_4, c_2_24_4;
    csa u_csa_2_24_4(s_1_24_8,s_1_24_7,s_1_24_6,s_2_24_4,c_2_24_4);
    wire s_2_24_5, c_2_24_5;
    csa u_csa_2_24_5(s_1_24_5,c_1_23_9,c_1_23_8,s_2_24_5,c_2_24_5);
    wire s_2_24_6, c_2_24_6;
    csa u_csa_2_24_6(c_1_23_7,c_1_23_6,c_1_23_5,s_2_24_6,c_2_24_6);
    wire s_2_25_4, c_2_25_4;
    csa u_csa_2_25_4(s_1_25_10,s_1_25_9,s_1_25_8,s_2_25_4,c_2_25_4);
    wire s_2_25_5, c_2_25_5;
    csa u_csa_2_25_5(s_1_25_7,s_1_25_6,s_1_25_5,s_2_25_5,c_2_25_5);
    wire s_2_25_6, c_2_25_6;
    csa u_csa_2_25_6(c_1_24_9,c_1_24_8,c_1_24_7,s_2_25_6,c_2_25_6);
    wire s_2_26_3, c_2_26_3;
    csa u_csa_2_26_3(c_0_25_8,c_0_25_9,s_1_26_10,s_2_26_3,c_2_26_3);
    wire s_2_26_4, c_2_26_4;
    csa u_csa_2_26_4(s_1_26_9,s_1_26_8,s_1_26_7,s_2_26_4,c_2_26_4);
    wire s_2_26_5, c_2_26_5;
    csa u_csa_2_26_5(s_1_26_6,c_1_25_10,c_1_25_9,s_2_26_5,c_2_26_5);
    wire s_2_26_6, c_2_26_6;
    csa u_csa_2_26_6(c_1_25_8,c_1_25_7,c_1_25_6,s_2_26_6,c_2_26_6);
    wire s_2_27_4, c_2_27_4;
    csa u_csa_2_27_4(c_0_26_8,s_1_27_9,s_1_27_8,s_2_27_4,c_2_27_4);
    wire s_2_27_5, c_2_27_5;
    csa u_csa_2_27_5(s_1_27_7,s_1_27_6,s_1_27_5,s_2_27_5,c_2_27_5);
    wire s_2_27_6, c_2_27_6;
    csa u_csa_2_27_6(c_1_26_10,c_1_26_9,c_1_26_8,s_2_27_6,c_2_27_6);
    wire s_2_28_3, c_2_28_3;
    csa u_csa_2_28_3(c_0_27_8,c_0_27_9,s_1_28_9,s_2_28_3,c_2_28_3);
    wire s_2_28_4, c_2_28_4;
    csa u_csa_2_28_4(s_1_28_8,s_1_28_7,s_1_28_6,s_2_28_4,c_2_28_4);
    wire s_2_28_5, c_2_28_5;
    csa u_csa_2_28_5(s_1_28_5,c_1_27_9,c_1_27_8,s_2_28_5,c_2_28_5);
    wire s_2_28_6, c_2_28_6;
    csa u_csa_2_28_6(c_1_27_7,c_1_27_6,c_1_27_5,s_2_28_6,c_2_28_6);
    wire s_2_29_4, c_2_29_4;
    csa u_csa_2_29_4(s_1_29_9,s_1_29_8,s_1_29_7,s_2_29_4,c_2_29_4);
    wire s_2_29_5, c_2_29_5;
    csa u_csa_2_29_5(s_1_29_6,s_1_29_5,c_1_28_9,s_2_29_5,c_2_29_5);
    wire s_2_29_6, c_2_29_6;
    csa u_csa_2_29_6(c_1_28_8,c_1_28_7,c_1_28_6,s_2_29_6,c_2_29_6);
    wire s_2_30_3, c_2_30_3;
    csa u_csa_2_30_3(c_0_29_7,c_0_29_8,s_1_30_8,s_2_30_3,c_2_30_3);
    wire s_2_30_4, c_2_30_4;
    csa u_csa_2_30_4(s_1_30_7,s_1_30_6,s_1_30_5,s_2_30_4,c_2_30_4);
    wire s_2_30_5, c_2_30_5;
    csa u_csa_2_30_5(c_1_29_9,c_1_29_8,c_1_29_7,s_2_30_5,c_2_30_5);
    wire s_2_31_3, c_2_31_3;
    csa u_csa_2_31_3(s_1_31_8,s_1_31_7,s_1_31_6,s_2_31_3,c_2_31_3);
    wire s_2_31_4, c_2_31_4;
    csa u_csa_2_31_4(s_1_31_5,s_1_31_4,c_1_30_8,s_2_31_4,c_2_31_4);
    wire s_2_31_5, c_2_31_5;
    csa u_csa_2_31_5(c_1_30_7,c_1_30_6,c_1_30_5,s_2_31_5,c_2_31_5);
    wire s_2_32_3, c_2_32_3;
    csa u_csa_2_32_3(c_0_31_7,s_1_32_8,s_1_32_7,s_2_32_3,c_2_32_3);
    wire s_2_32_4, c_2_32_4;
    csa u_csa_2_32_4(s_1_32_6,s_1_32_5,c_1_31_8,s_2_32_4,c_2_32_4);
    wire s_2_32_5, c_2_32_5;
    csa u_csa_2_32_5(c_1_31_7,c_1_31_6,c_1_31_5,s_2_32_5,c_2_32_5);
    wire s_2_33_3, c_2_33_3;
    csa u_csa_2_33_3(s_1_33_7,s_1_33_6,s_1_33_5,s_2_33_3,c_2_33_3);
    wire s_2_33_4, c_2_33_4;
    csa u_csa_2_33_4(s_1_33_4,c_1_32_8,c_1_32_7,s_2_33_4,c_2_33_4);
    wire s_2_34_2, c_2_34_2;
    csa u_csa_2_34_2(c_0_33_6,s_1_34_7,s_1_34_6,s_2_34_2,c_2_34_2);
    wire s_2_34_3, c_2_34_3;
    csa u_csa_2_34_3(s_1_34_5,s_1_34_4,c_1_33_7,s_2_34_3,c_2_34_3);
    wire s_2_34_4, c_2_34_4;
    csa u_csa_2_34_4(c_1_33_6,c_1_33_5,c_1_33_4,s_2_34_4,c_2_34_4);
    wire s_2_35_3, c_2_35_3;
    csa u_csa_2_35_3(c_0_34_6,c_0_34_7,s_1_35_6,s_2_35_3,c_2_35_3);
    wire s_2_35_4, c_2_35_4;
    csa u_csa_2_35_4(s_1_35_5,s_1_35_4,c_1_34_7,s_2_35_4,c_2_35_4);
    wire s_2_35_5, c_2_35_5;
    csa u_csa_2_35_5(c_1_34_6,c_1_34_5,c_1_34_4,s_2_35_5,c_2_35_5);
    wire s_2_36_3, c_2_36_3;
    csa u_csa_2_36_3(c_0_35_5,s_1_36_5,s_1_36_4,s_2_36_3,c_2_36_3);
    wire s_2_36_4, c_2_36_4;
    csa u_csa_2_36_4(s_1_36_3,c_1_35_6,c_1_35_5,s_2_36_4,c_2_36_4);
    wire s_2_37_2, c_2_37_2;
    csa u_csa_2_37_2(c_0_36_5,c_0_36_6,s_1_37_5,s_2_37_2,c_2_37_2);
    wire s_2_37_3, c_2_37_3;
    csa u_csa_2_37_3(s_1_37_4,s_1_37_3,c_1_36_5,s_2_37_3,c_2_37_3);
    wire s_2_38_2, c_2_38_2;
    csa u_csa_2_38_2(s_1_38_5,s_1_38_4,s_1_38_3,s_2_38_2,c_2_38_2);
    wire s_2_38_3, c_2_38_3;
    csa u_csa_2_38_3(c_1_37_5,c_1_37_4,c_1_37_3,s_2_38_3,c_2_38_3);
    wire s_2_39_2, c_2_39_2;
    csa u_csa_2_39_2(c_0_38_4,c_0_38_5,s_1_39_4,s_2_39_2,c_2_39_2);
    wire s_2_39_3, c_2_39_3;
    csa u_csa_2_39_3(s_1_39_3,c_1_38_5,c_1_38_4,s_2_39_3,c_2_39_3);
    wire s_2_40_2, c_2_40_2;
    csa u_csa_2_40_2(s_1_40_4,s_1_40_3,s_1_40_2,s_2_40_2,c_2_40_2);
    wire s_2_41_1, c_2_41_1;
    csa u_csa_2_41_1(c_0_40_4,s_1_41_4,s_1_41_3,s_2_41_1,c_2_41_1);
    wire s_2_41_2, c_2_41_2;
    csa u_csa_2_41_2(c_1_40_4,c_1_40_3,c_1_40_2,s_2_41_2,c_2_41_2);
    wire s_2_42_2, c_2_42_2;
    csa u_csa_2_42_2(s_1_42_3,s_1_42_2,c_1_41_4,s_2_42_2,c_2_42_2);
    wire s_2_43_1, c_2_43_1;
    csa u_csa_2_43_1(c_0_42_3,s_1_43_3,s_1_43_2,s_2_43_1,c_2_43_1);
    wire s_2_44_1, c_2_44_1;
    csa u_csa_2_44_1(c_0_43_3,c_0_43_4,s_1_44_2,s_2_44_1,c_2_44_1);
    wire s_2_45_1, c_2_45_1;
    csa u_csa_2_45_1(c_0_44_2,s_1_45_1,c_1_44_2,s_2_45_1,c_2_45_1);
    wire s_2_46_1, c_2_46_1;
    csa u_csa_2_46_1(c_0_45_2,c_0_45_3,s_1_46_1,s_2_46_1,c_2_46_1);
    wire s_2_48_0, c_2_48_0;
    csa u_csa_2_48_0(c_0_47_1,s_0_48_1,c_1_47_1,s_2_48_0,c_2_48_0);
    wire s_3_5_0, c_3_5_0;
    csa u_csa_3_5_0(c_1_4_1,s_1_5_1,c_2_4_0,s_3_5_0,c_3_5_0);
    wire s_3_8_0, c_3_8_0;
    csa u_csa_3_8_0(c_1_7_1,c_1_7_2,s_2_8_1,s_3_8_0,c_3_8_0);
    wire s_3_9_1, c_3_9_1;
    csa u_csa_3_9_1(c_1_8_2,s_2_9_1,c_2_8_1,s_3_9_1,c_3_9_1);
    wire s_3_10_1, c_3_10_1;
    csa u_csa_3_10_1(s_2_10_2,s_2_10_1,c_2_9_1,s_3_10_1,c_3_10_1);
    wire s_3_11_1, c_3_11_1;
    csa u_csa_3_11_1(c_1_10_2,c_1_10_3,s_2_11_2,s_3_11_1,c_3_11_1);
    wire s_3_12_1, c_3_12_1;
    csa u_csa_3_12_1(c_1_11_2,c_1_11_3,s_2_12_1,s_3_12_1,c_3_12_1);
    wire s_3_13_1, c_3_13_1;
    csa u_csa_3_13_1(c_1_12_2,s_2_13_2,s_2_13_1,s_3_13_1,c_3_13_1);
    wire s_3_14_1, c_3_14_1;
    csa u_csa_3_14_1(s_2_14_3,s_2_14_2,c_2_13_2,s_3_14_1,c_3_14_1);
    wire s_3_15_1, c_3_15_1;
    csa u_csa_3_15_1(c_1_14_3,c_1_14_4,s_2_15_3,s_3_15_1,c_3_15_1);
    wire s_3_15_2, c_3_15_2;
    csa u_csa_3_15_2(s_2_15_2,c_2_14_3,c_2_14_2,s_3_15_2,c_3_15_2);
    wire s_3_16_2, c_3_16_2;
    csa u_csa_3_16_2(c_1_15_3,s_2_16_3,s_2_16_2,s_3_16_2,c_3_16_2);
    wire s_3_17_1, c_3_17_1;
    csa u_csa_3_17_1(s_2_17_4,s_2_17_3,s_2_17_2,s_3_17_1,c_3_17_1);
    wire s_3_18_1, c_3_18_1;
    csa u_csa_3_18_1(c_1_17_4,c_1_17_5,s_2_18_4,s_3_18_1,c_3_18_1);
    wire s_3_18_2, c_3_18_2;
    csa u_csa_3_18_2(s_2_18_3,c_2_17_4,c_2_17_3,s_3_18_2,c_3_18_2);
    wire s_3_19_2, c_3_19_2;
    csa u_csa_3_19_2(c_1_18_3,s_2_19_4,s_2_19_3,s_3_19_2,c_3_19_2);
    wire s_3_19_3, c_3_19_3;
    csa u_csa_3_19_3(s_2_19_2,c_2_18_4,c_2_18_3,s_3_19_3,c_3_19_3);
    wire s_3_20_2, c_3_20_2;
    csa u_csa_3_20_2(s_2_20_5,s_2_20_4,s_2_20_3,s_3_20_2,c_3_20_2);
    wire s_3_20_3, c_3_20_3;
    csa u_csa_3_20_3(c_2_19_4,c_2_19_3,c_2_19_2,s_3_20_3,c_3_20_3);
    wire s_3_21_2, c_3_21_2;
    csa u_csa_3_21_2(s_2_21_5,s_2_21_4,s_2_21_3,s_3_21_2,c_3_21_2);
    wire s_3_21_3, c_3_21_3;
    csa u_csa_3_21_3(c_2_20_5,c_2_20_4,c_2_20_3,s_3_21_3,c_3_21_3);
    wire s_3_22_2, c_3_22_2;
    csa u_csa_3_22_2(c_1_21_4,c_1_21_5,s_2_22_5,s_3_22_2,c_3_22_2);
    wire s_3_22_3, c_3_22_3;
    csa u_csa_3_22_3(s_2_22_4,s_2_22_3,c_2_21_5,s_3_22_3,c_3_22_3);
    wire s_3_23_2, c_3_23_2;
    csa u_csa_3_23_2(c_1_22_5,s_2_23_5,s_2_23_4,s_3_23_2,c_3_23_2);
    wire s_3_23_3, c_3_23_3;
    csa u_csa_3_23_3(s_2_23_3,c_2_22_5,c_2_22_4,s_3_23_3,c_3_23_3);
    wire s_3_24_2, c_3_24_2;
    csa u_csa_3_24_2(s_2_24_6,s_2_24_5,s_2_24_4,s_3_24_2,c_3_24_2);
    wire s_3_24_3, c_3_24_3;
    csa u_csa_3_24_3(s_2_24_3,c_2_23_5,c_2_23_4,s_3_24_3,c_3_24_3);
    wire s_3_25_2, c_3_25_2;
    csa u_csa_3_25_2(c_1_24_5,c_1_24_6,s_2_25_6,s_3_25_2,c_3_25_2);
    wire s_3_25_3, c_3_25_3;
    csa u_csa_3_25_3(s_2_25_5,s_2_25_4,c_2_24_6,s_3_25_3,c_3_25_3);
    wire s_3_25_4, c_3_25_4;
    csa u_csa_3_25_4(c_2_24_5,c_2_24_4,c_2_24_3,s_3_25_4,c_3_25_4);
    wire s_3_26_3, c_3_26_3;
    csa u_csa_3_26_3(c_1_25_5,s_2_26_6,s_2_26_5,s_3_26_3,c_3_26_3);
    wire s_3_26_4, c_3_26_4;
    csa u_csa_3_26_4(s_2_26_4,s_2_26_3,c_2_25_6,s_3_26_4,c_3_26_4);
    wire s_3_27_2, c_3_27_2;
    csa u_csa_3_27_2(c_1_26_6,c_1_26_7,s_2_27_6,s_3_27_2,c_3_27_2);
    wire s_3_27_3, c_3_27_3;
    csa u_csa_3_27_3(s_2_27_5,s_2_27_4,c_2_26_6,s_3_27_3,c_3_27_3);
    wire s_3_27_4, c_3_27_4;
    csa u_csa_3_27_4(c_2_26_5,c_2_26_4,c_2_26_3,s_3_27_4,c_3_27_4);
    wire s_3_28_3, c_3_28_3;
    csa u_csa_3_28_3(s_2_28_6,s_2_28_5,s_2_28_4,s_3_28_3,c_3_28_3);
    wire s_3_28_4, c_3_28_4;
    csa u_csa_3_28_4(s_2_28_3,c_2_27_6,c_2_27_5,s_3_28_4,c_3_28_4);
    wire s_3_29_2, c_3_29_2;
    csa u_csa_3_29_2(c_1_28_5,s_2_29_6,s_2_29_5,s_3_29_2,c_3_29_2);
    wire s_3_29_3, c_3_29_3;
    csa u_csa_3_29_3(s_2_29_4,c_2_28_6,c_2_28_5,s_3_29_3,c_3_29_3);
    wire s_3_30_2, c_3_30_2;
    csa u_csa_3_30_2(c_1_29_5,c_1_29_6,s_2_30_5,s_3_30_2,c_3_30_2);
    wire s_3_30_3, c_3_30_3;
    csa u_csa_3_30_3(s_2_30_4,s_2_30_3,c_2_29_6,s_3_30_3,c_3_30_3);
    wire s_3_31_2, c_3_31_2;
    csa u_csa_3_31_2(s_2_31_5,s_2_31_4,s_2_31_3,s_3_31_2,c_3_31_2);
    wire s_3_31_3, c_3_31_3;
    csa u_csa_3_31_3(c_2_30_5,c_2_30_4,c_2_30_3,s_3_31_3,c_3_31_3);
    wire s_3_32_2, c_3_32_2;
    csa u_csa_3_32_2(c_1_31_4,s_2_32_5,s_2_32_4,s_3_32_2,c_3_32_2);
    wire s_3_32_3, c_3_32_3;
    csa u_csa_3_32_3(s_2_32_3,c_2_31_5,c_2_31_4,s_3_32_3,c_3_32_3);
    wire s_3_33_2, c_3_33_2;
    csa u_csa_3_33_2(c_1_32_5,c_1_32_6,s_2_33_4,s_3_33_2,c_3_33_2);
    wire s_3_33_3, c_3_33_3;
    csa u_csa_3_33_3(s_2_33_3,c_2_32_5,c_2_32_4,s_3_33_3,c_3_33_3);
    wire s_3_34_2, c_3_34_2;
    csa u_csa_3_34_2(s_2_34_4,s_2_34_3,s_2_34_2,s_3_34_2,c_3_34_2);
    wire s_3_35_1, c_3_35_1;
    csa u_csa_3_35_1(s_2_35_5,s_2_35_4,s_2_35_3,s_3_35_1,c_3_35_1);
    wire s_3_35_2, c_3_35_2;
    csa u_csa_3_35_2(c_2_34_4,c_2_34_3,c_2_34_2,s_3_35_2,c_3_35_2);
    wire s_3_36_2, c_3_36_2;
    csa u_csa_3_36_2(c_1_35_4,s_2_36_4,s_2_36_3,s_3_36_2,c_3_36_2);
    wire s_3_36_3, c_3_36_3;
    csa u_csa_3_36_3(c_2_35_5,c_2_35_4,c_2_35_3,s_3_36_3,c_3_36_3);
    wire s_3_37_2, c_3_37_2;
    csa u_csa_3_37_2(c_1_36_3,c_1_36_4,s_2_37_3,s_3_37_2,c_3_37_2);
    wire s_3_37_3, c_3_37_3;
    csa u_csa_3_37_3(s_2_37_2,c_2_36_4,c_2_36_3,s_3_37_3,c_3_37_3);
    wire s_3_38_2, c_3_38_2;
    csa u_csa_3_38_2(s_2_38_3,s_2_38_2,c_2_37_3,s_3_38_2,c_3_38_2);
    wire s_3_39_1, c_3_39_1;
    csa u_csa_3_39_1(c_1_38_3,s_2_39_3,s_2_39_2,s_3_39_1,c_3_39_1);
    wire s_3_40_1, c_3_40_1;
    csa u_csa_3_40_1(c_1_39_3,c_1_39_4,s_2_40_2,s_3_40_1,c_3_40_1);
    wire s_3_41_1, c_3_41_1;
    csa u_csa_3_41_1(s_2_41_2,s_2_41_1,c_2_40_2,s_3_41_1,c_3_41_1);
    wire s_3_42_1, c_3_42_1;
    csa u_csa_3_42_1(c_1_41_3,s_2_42_2,c_2_41_2,s_3_42_1,c_3_42_1);
    wire s_3_43_1, c_3_43_1;
    csa u_csa_3_43_1(c_1_42_2,c_1_42_3,s_2_43_1,s_3_43_1,c_3_43_1);
    wire s_3_44_1, c_3_44_1;
    csa u_csa_3_44_1(c_1_43_2,c_1_43_3,s_2_44_1,s_3_44_1,c_3_44_1);
    wire s_3_46_0, c_3_46_0;
    csa u_csa_3_46_0(c_1_45_1,s_2_46_1,c_2_45_1,s_3_46_0,c_3_46_0);
    wire s_3_47_1, c_3_47_1;
    csa u_csa_3_47_1(c_1_46_1,s_1_47_1,c_2_46_1,s_3_47_1,c_3_47_1);
    wire s_4_6_0, c_4_6_0;
    csa u_csa_4_6_0(s_2_6_0,c_1_5_1,c_3_5_0,s_4_6_0,c_4_6_0);
    wire s_4_11_0, c_4_11_0;
    csa u_csa_4_11_0(c_2_10_1,c_2_10_2,s_3_11_1,s_4_11_0,c_4_11_0);
    wire s_4_12_1, c_4_12_1;
    csa u_csa_4_12_1(c_2_11_2,s_3_12_1,c_3_11_1,s_4_12_1,c_4_12_1);
    wire s_4_13_1, c_4_13_1;
    csa u_csa_4_13_1(c_2_12_1,s_3_13_1,c_3_12_1,s_4_13_1,c_4_13_1);
    wire s_4_14_1, c_4_14_1;
    csa u_csa_4_14_1(c_2_13_1,s_3_14_1,c_3_13_1,s_4_14_1,c_4_14_1);
    wire s_4_15_1, c_4_15_1;
    csa u_csa_4_15_1(s_3_15_2,s_3_15_1,c_3_14_1,s_4_15_1,c_4_15_1);
    wire s_4_16_1, c_4_16_1;
    csa u_csa_4_16_1(c_2_15_2,c_2_15_3,s_3_16_2,s_4_16_1,c_4_16_1);
    wire s_4_17_1, c_4_17_1;
    csa u_csa_4_17_1(c_2_16_2,c_2_16_3,s_3_17_1,s_4_17_1,c_4_17_1);
    wire s_4_18_1, c_4_18_1;
    csa u_csa_4_18_1(c_2_17_2,s_3_18_2,s_3_18_1,s_4_18_1,c_4_18_1);
    wire s_4_19_1, c_4_19_1;
    csa u_csa_4_19_1(s_3_19_3,s_3_19_2,c_3_18_2,s_4_19_1,c_4_19_1);
    wire s_4_20_1, c_4_20_1;
    csa u_csa_4_20_1(s_3_20_3,s_3_20_2,c_3_19_3,s_4_20_1,c_4_20_1);
    wire s_4_21_1, c_4_21_1;
    csa u_csa_4_21_1(s_3_21_3,s_3_21_2,c_3_20_3,s_4_21_1,c_4_21_1);
    wire s_4_22_1, c_4_22_1;
    csa u_csa_4_22_1(c_2_21_3,c_2_21_4,s_3_22_3,s_4_22_1,c_4_22_1);
    wire s_4_22_2, c_4_22_2;
    csa u_csa_4_22_2(s_3_22_2,c_3_21_3,c_3_21_2,s_4_22_2,c_4_22_2);
    wire s_4_23_2, c_4_23_2;
    csa u_csa_4_23_2(c_2_22_3,s_3_23_3,s_3_23_2,s_4_23_2,c_4_23_2);
    wire s_4_24_1, c_4_24_1;
    csa u_csa_4_24_1(c_2_23_3,s_3_24_3,s_3_24_2,s_4_24_1,c_4_24_1);
    wire s_4_25_1, c_4_25_1;
    csa u_csa_4_25_1(s_3_25_4,s_3_25_3,s_3_25_2,s_4_25_1,c_4_25_1);
    wire s_4_26_1, c_4_26_1;
    csa u_csa_4_26_1(c_2_25_4,c_2_25_5,s_3_26_4,s_4_26_1,c_4_26_1);
    wire s_4_26_2, c_4_26_2;
    csa u_csa_4_26_2(s_3_26_3,c_3_25_4,c_3_25_3,s_4_26_2,c_4_26_2);
    wire s_4_27_2, c_4_27_2;
    csa u_csa_4_27_2(s_3_27_4,s_3_27_3,s_3_27_2,s_4_27_2,c_4_27_2);
    wire s_4_28_1, c_4_28_1;
    csa u_csa_4_28_1(c_2_27_4,s_3_28_4,s_3_28_3,s_4_28_1,c_4_28_1);
    wire s_4_28_2, c_4_28_2;
    csa u_csa_4_28_2(c_3_27_4,c_3_27_3,c_3_27_2,s_4_28_2,c_4_28_2);
    wire s_4_29_2, c_4_29_2;
    csa u_csa_4_29_2(c_2_28_3,c_2_28_4,s_3_29_3,s_4_29_2,c_4_29_2);
    wire s_4_29_3, c_4_29_3;
    csa u_csa_4_29_3(s_3_29_2,c_3_28_4,c_3_28_3,s_4_29_3,c_4_29_3);
    wire s_4_30_2, c_4_30_2;
    csa u_csa_4_30_2(c_2_29_4,c_2_29_5,s_3_30_3,s_4_30_2,c_4_30_2);
    wire s_4_30_3, c_4_30_3;
    csa u_csa_4_30_3(s_3_30_2,c_3_29_3,c_3_29_2,s_4_30_3,c_4_30_3);
    wire s_4_31_2, c_4_31_2;
    csa u_csa_4_31_2(s_3_31_3,s_3_31_2,c_3_30_3,s_4_31_2,c_4_31_2);
    wire s_4_32_1, c_4_32_1;
    csa u_csa_4_32_1(c_2_31_3,s_3_32_3,s_3_32_2,s_4_32_1,c_4_32_1);
    wire s_4_33_1, c_4_33_1;
    csa u_csa_4_33_1(c_2_32_3,s_3_33_3,s_3_33_2,s_4_33_1,c_4_33_1);
    wire s_4_34_1, c_4_34_1;
    csa u_csa_4_34_1(c_2_33_3,c_2_33_4,s_3_34_2,s_4_34_1,c_4_34_1);
    wire s_4_35_1, c_4_35_1;
    csa u_csa_4_35_1(s_3_35_2,s_3_35_1,c_3_34_2,s_4_35_1,c_4_35_1);
    wire s_4_36_1, c_4_36_1;
    csa u_csa_4_36_1(s_3_36_3,s_3_36_2,c_3_35_2,s_4_36_1,c_4_36_1);
    wire s_4_37_1, c_4_37_1;
    csa u_csa_4_37_1(s_3_37_3,s_3_37_2,c_3_36_3,s_4_37_1,c_4_37_1);
    wire s_4_38_1, c_4_38_1;
    csa u_csa_4_38_1(c_2_37_2,s_3_38_2,c_3_37_3,s_4_38_1,c_4_38_1);
    wire s_4_39_1, c_4_39_1;
    csa u_csa_4_39_1(c_2_38_2,c_2_38_3,s_3_39_1,s_4_39_1,c_4_39_1);
    wire s_4_40_1, c_4_40_1;
    csa u_csa_4_40_1(c_2_39_2,c_2_39_3,s_3_40_1,s_4_40_1,c_4_40_1);
    wire s_4_42_0, c_4_42_0;
    csa u_csa_4_42_0(c_2_41_1,s_3_42_1,c_3_41_1,s_4_42_0,c_4_42_0);
    wire s_4_43_1, c_4_43_1;
    csa u_csa_4_43_1(c_2_42_2,s_3_43_1,c_3_42_1,s_4_43_1,c_4_43_1);
    wire s_4_44_1, c_4_44_1;
    csa u_csa_4_44_1(c_2_43_1,s_3_44_1,c_3_43_1,s_4_44_1,c_4_44_1);
    wire s_4_45_1, c_4_45_1;
    csa u_csa_4_45_1(c_2_44_1,s_2_45_1,c_3_44_1,s_4_45_1,c_4_45_1);
    wire s_5_7_0, c_5_7_0;
    csa u_csa_5_7_0(s_2_7_1,c_2_6_0,c_4_6_0,s_5_7_0,c_5_7_0);
    wire s_5_16_0, c_5_16_0;
    csa u_csa_5_16_0(c_3_15_1,c_3_15_2,s_4_16_1,s_5_16_0,c_5_16_0);
    wire s_5_17_1, c_5_17_1;
    csa u_csa_5_17_1(c_3_16_2,s_4_17_1,c_4_16_1,s_5_17_1,c_5_17_1);
    wire s_5_18_1, c_5_18_1;
    csa u_csa_5_18_1(c_3_17_1,s_4_18_1,c_4_17_1,s_5_18_1,c_5_18_1);
    wire s_5_19_1, c_5_19_1;
    csa u_csa_5_19_1(c_3_18_1,s_4_19_1,c_4_18_1,s_5_19_1,c_5_19_1);
    wire s_5_20_1, c_5_20_1;
    csa u_csa_5_20_1(c_3_19_2,s_4_20_1,c_4_19_1,s_5_20_1,c_5_20_1);
    wire s_5_21_1, c_5_21_1;
    csa u_csa_5_21_1(c_3_20_2,s_4_21_1,c_4_20_1,s_5_21_1,c_5_21_1);
    wire s_5_22_1, c_5_22_1;
    csa u_csa_5_22_1(s_4_22_2,s_4_22_1,c_4_21_1,s_5_22_1,c_5_22_1);
    wire s_5_23_1, c_5_23_1;
    csa u_csa_5_23_1(c_3_22_2,c_3_22_3,s_4_23_2,s_5_23_1,c_5_23_1);
    wire s_5_24_1, c_5_24_1;
    csa u_csa_5_24_1(c_3_23_2,c_3_23_3,s_4_24_1,s_5_24_1,c_5_24_1);
    wire s_5_25_1, c_5_25_1;
    csa u_csa_5_25_1(c_3_24_2,c_3_24_3,s_4_25_1,s_5_25_1,c_5_25_1);
    wire s_5_26_1, c_5_26_1;
    csa u_csa_5_26_1(c_3_25_2,s_4_26_2,s_4_26_1,s_5_26_1,c_5_26_1);
    wire s_5_27_1, c_5_27_1;
    csa u_csa_5_27_1(c_3_26_3,c_3_26_4,s_4_27_2,s_5_27_1,c_5_27_1);
    wire s_5_28_1, c_5_28_1;
    csa u_csa_5_28_1(s_4_28_2,s_4_28_1,c_4_27_2,s_5_28_1,c_5_28_1);
    wire s_5_29_1, c_5_29_1;
    csa u_csa_5_29_1(s_4_29_3,s_4_29_2,c_4_28_2,s_5_29_1,c_5_29_1);
    wire s_5_30_1, c_5_30_1;
    csa u_csa_5_30_1(s_4_30_3,s_4_30_2,c_4_29_3,s_5_30_1,c_5_30_1);
    wire s_5_31_1, c_5_31_1;
    csa u_csa_5_31_1(c_3_30_2,s_4_31_2,c_4_30_3,s_5_31_1,c_5_31_1);
    wire s_5_32_1, c_5_32_1;
    csa u_csa_5_32_1(c_3_31_2,c_3_31_3,s_4_32_1,s_5_32_1,c_5_32_1);
    wire s_5_33_1, c_5_33_1;
    csa u_csa_5_33_1(c_3_32_2,c_3_32_3,s_4_33_1,s_5_33_1,c_5_33_1);
    wire s_5_34_1, c_5_34_1;
    csa u_csa_5_34_1(c_3_33_2,c_3_33_3,s_4_34_1,s_5_34_1,c_5_34_1);
    wire s_5_36_0, c_5_36_0;
    csa u_csa_5_36_0(c_3_35_1,s_4_36_1,c_4_35_1,s_5_36_0,c_5_36_0);
    wire s_5_37_1, c_5_37_1;
    csa u_csa_5_37_1(c_3_36_2,s_4_37_1,c_4_36_1,s_5_37_1,c_5_37_1);
    wire s_5_38_1, c_5_38_1;
    csa u_csa_5_38_1(c_3_37_2,s_4_38_1,c_4_37_1,s_5_38_1,c_5_38_1);
    wire s_5_39_1, c_5_39_1;
    csa u_csa_5_39_1(c_3_38_2,s_4_39_1,c_4_38_1,s_5_39_1,c_5_39_1);
    wire s_5_40_1, c_5_40_1;
    csa u_csa_5_40_1(c_3_39_1,s_4_40_1,c_4_39_1,s_5_40_1,c_5_40_1);
    wire s_5_41_1, c_5_41_1;
    csa u_csa_5_41_1(c_3_40_1,s_3_41_1,c_4_40_1,s_5_41_1,c_5_41_1);
    wire s_6_8_0, c_6_8_0;
    csa u_csa_6_8_0(c_2_7_1,s_3_8_0,c_5_7_0,s_6_8_0,c_6_8_0);
    wire s_6_23_0, c_6_23_0;
    csa u_csa_6_23_0(c_4_22_1,c_4_22_2,s_5_23_1,s_6_23_0,c_6_23_0);
    wire s_6_24_1, c_6_24_1;
    csa u_csa_6_24_1(c_4_23_2,s_5_24_1,c_5_23_1,s_6_24_1,c_6_24_1);
    wire s_6_25_1, c_6_25_1;
    csa u_csa_6_25_1(c_4_24_1,s_5_25_1,c_5_24_1,s_6_25_1,c_6_25_1);
    wire s_6_26_1, c_6_26_1;
    csa u_csa_6_26_1(c_4_25_1,s_5_26_1,c_5_25_1,s_6_26_1,c_6_26_1);
    wire s_6_27_1, c_6_27_1;
    csa u_csa_6_27_1(c_4_26_1,c_4_26_2,s_5_27_1,s_6_27_1,c_6_27_1);
    wire s_6_29_0, c_6_29_0;
    csa u_csa_6_29_0(c_4_28_1,s_5_29_1,c_5_28_1,s_6_29_0,c_6_29_0);
    wire s_6_30_1, c_6_30_1;
    csa u_csa_6_30_1(c_4_29_2,s_5_30_1,c_5_29_1,s_6_30_1,c_6_30_1);
    wire s_6_31_1, c_6_31_1;
    csa u_csa_6_31_1(c_4_30_2,s_5_31_1,c_5_30_1,s_6_31_1,c_6_31_1);
    wire s_6_32_1, c_6_32_1;
    csa u_csa_6_32_1(c_4_31_2,s_5_32_1,c_5_31_1,s_6_32_1,c_6_32_1);
    wire s_6_33_1, c_6_33_1;
    csa u_csa_6_33_1(c_4_32_1,s_5_33_1,c_5_32_1,s_6_33_1,c_6_33_1);
    wire s_6_34_1, c_6_34_1;
    csa u_csa_6_34_1(c_4_33_1,s_5_34_1,c_5_33_1,s_6_34_1,c_6_34_1);
    wire s_6_35_1, c_6_35_1;
    csa u_csa_6_35_1(c_4_34_1,s_4_35_1,c_5_34_1,s_6_35_1,c_6_35_1);
    wire s_7_9_0, c_7_9_0;
    csa u_csa_7_9_0(c_3_8_0,s_3_9_1,c_6_8_0,s_7_9_0,c_7_9_0);
    wire s_7_27_0, c_7_27_0;
    csa u_csa_7_27_0(c_5_26_1,s_6_27_1,c_6_26_1,s_7_27_0,c_7_27_0);
    wire s_7_28_1, c_7_28_1;
    csa u_csa_7_28_1(c_5_27_1,s_5_28_1,c_6_27_1,s_7_28_1,c_7_28_1);
    wire s_8_10_0, c_8_10_0;
    csa u_csa_8_10_0(s_3_10_1,c_3_9_1,c_7_9_0,s_8_10_0,c_8_10_0);
    wire s_9_11_0, c_9_11_0;
    csa u_csa_9_11_0(c_3_10_1,s_4_11_0,c_8_10_0,s_9_11_0,c_9_11_0);
    wire s_10_12_0, c_10_12_0;
    csa u_csa_10_12_0(c_4_11_0,s_4_12_1,c_9_11_0,s_10_12_0,c_10_12_0);
    wire s_11_13_0, c_11_13_0;
    csa u_csa_11_13_0(s_4_13_1,c_4_12_1,c_10_12_0,s_11_13_0,c_11_13_0);
    wire s_12_14_0, c_12_14_0;
    csa u_csa_12_14_0(c_4_13_1,s_4_14_1,c_11_13_0,s_12_14_0,c_12_14_0);
    wire s_13_15_0, c_13_15_0;
    csa u_csa_13_15_0(s_4_15_1,c_4_14_1,c_12_14_0,s_13_15_0,c_13_15_0);
    wire s_14_16_0, c_14_16_0;
    csa u_csa_14_16_0(c_4_15_1,s_5_16_0,c_13_15_0,s_14_16_0,c_14_16_0);
    wire s_15_17_0, c_15_17_0;
    csa u_csa_15_17_0(c_5_16_0,s_5_17_1,c_14_16_0,s_15_17_0,c_15_17_0);
    wire s_16_18_0, c_16_18_0;
    csa u_csa_16_18_0(s_5_18_1,c_5_17_1,c_15_17_0,s_16_18_0,c_16_18_0);
    wire s_17_19_0, c_17_19_0;
    csa u_csa_17_19_0(c_5_18_1,s_5_19_1,c_16_18_0,s_17_19_0,c_17_19_0);
    wire s_18_20_0, c_18_20_0;
    csa u_csa_18_20_0(s_5_20_1,c_5_19_1,c_17_19_0,s_18_20_0,c_18_20_0);
    wire s_19_21_0, c_19_21_0;
    csa u_csa_19_21_0(c_5_20_1,s_5_21_1,c_18_20_0,s_19_21_0,c_19_21_0);
    wire s_20_22_0, c_20_22_0;
    csa u_csa_20_22_0(s_5_22_1,c_5_21_1,c_19_21_0,s_20_22_0,c_20_22_0);
    wire s_21_23_0, c_21_23_0;
    csa u_csa_21_23_0(c_5_22_1,s_6_23_0,c_20_22_0,s_21_23_0,c_21_23_0);
    wire s_22_24_0, c_22_24_0;
    csa u_csa_22_24_0(c_6_23_0,s_6_24_1,c_21_23_0,s_22_24_0,c_22_24_0);
    wire s_23_25_0, c_23_25_0;
    csa u_csa_23_25_0(s_6_25_1,c_6_24_1,c_22_24_0,s_23_25_0,c_23_25_0);
    wire s_24_26_0, c_24_26_0;
    csa u_csa_24_26_0(c_6_25_1,s_6_26_1,c_23_25_0,s_24_26_0,c_24_26_0);

    wire [51:0] row0_vec;
    wire [51:0] row1_vec;
    assign row0_vec[0] = pp[0][0];
    assign row0_vec[1] = pp[0][1];
    assign row0_vec[2] = s_0_2_0;
    assign row0_vec[3] = s_1_3_0;
    assign row0_vec[4] = s_2_4_0;
    assign row0_vec[5] = s_3_5_0;
    assign row0_vec[6] = s_4_6_0;
    assign row0_vec[7] = s_5_7_0;
    assign row0_vec[8] = s_6_8_0;
    assign row0_vec[9] = s_7_9_0;
    assign row0_vec[10] = s_8_10_0;
    assign row0_vec[11] = s_9_11_0;
    assign row0_vec[12] = s_10_12_0;
    assign row0_vec[13] = s_11_13_0;
    assign row0_vec[14] = s_12_14_0;
    assign row0_vec[15] = s_13_15_0;
    assign row0_vec[16] = s_14_16_0;
    assign row0_vec[17] = s_15_17_0;
    assign row0_vec[18] = s_16_18_0;
    assign row0_vec[19] = s_17_19_0;
    assign row0_vec[20] = s_18_20_0;
    assign row0_vec[21] = s_19_21_0;
    assign row0_vec[22] = s_20_22_0;
    assign row0_vec[23] = s_21_23_0;
    assign row0_vec[24] = s_22_24_0;
    assign row0_vec[25] = s_23_25_0;
    assign row0_vec[26] = s_24_26_0;
    assign row0_vec[27] = s_7_27_0;
    assign row0_vec[28] = c_7_27_0;
    assign row0_vec[29] = c_7_28_1;
    assign row0_vec[30] = s_6_30_1;
    assign row0_vec[31] = s_6_31_1;
    assign row0_vec[32] = s_6_32_1;
    assign row0_vec[33] = s_6_33_1;
    assign row0_vec[34] = s_6_34_1;
    assign row0_vec[35] = s_6_35_1;
    assign row0_vec[36] = s_5_36_0;
    assign row0_vec[37] = c_5_36_0;
    assign row0_vec[38] = c_5_37_1;
    assign row0_vec[39] = c_5_38_1;
    assign row0_vec[40] = c_5_39_1;
    assign row0_vec[41] = c_5_40_1;
    assign row0_vec[42] = c_5_41_1;
    assign row0_vec[43] = s_4_43_1;
    assign row0_vec[44] = s_4_44_1;
    assign row0_vec[45] = s_4_45_1;
    assign row0_vec[46] = s_3_46_0;
    assign row0_vec[47] = c_3_46_0;
    assign row0_vec[48] = c_3_47_1;
    assign row0_vec[49] = s_1_49_0;
    assign row0_vec[50] = c_1_49_0;
    assign row0_vec[51] = 1'b0;
    assign row1_vec[1] = pp[1][0];
    assign row1_vec[27] = c_24_26_0;
    assign row1_vec[28] = s_7_28_1;
    assign row1_vec[29] = s_6_29_0;
    assign row1_vec[30] = c_6_29_0;
    assign row1_vec[31] = c_6_30_1;
    assign row1_vec[32] = c_6_31_1;
    assign row1_vec[33] = c_6_32_1;
    assign row1_vec[34] = c_6_33_1;
    assign row1_vec[35] = c_6_34_1;
    assign row1_vec[36] = c_6_35_1;
    assign row1_vec[37] = s_5_37_1;
    assign row1_vec[38] = s_5_38_1;
    assign row1_vec[39] = s_5_39_1;
    assign row1_vec[40] = s_5_40_1;
    assign row1_vec[41] = s_5_41_1;
    assign row1_vec[42] = s_4_42_0;
    assign row1_vec[43] = c_4_42_0;
    assign row1_vec[44] = c_4_43_1;
    assign row1_vec[45] = c_4_44_1;
    assign row1_vec[46] = c_4_45_1;
    assign row1_vec[47] = s_3_47_1;
    assign row1_vec[48] = s_2_48_0;
    assign row1_vec[49] = c_2_48_0;
    assign row1_vec[50] = pp[25][25];
    assign row1_vec[0] = 1'b0;
    assign row1_vec[2] = 1'b0;
    assign row1_vec[3] = 1'b0;
    assign row1_vec[4] = 1'b0;
    assign row1_vec[5] = 1'b0;
    assign row1_vec[6] = 1'b0;
    assign row1_vec[7] = 1'b0;
    assign row1_vec[8] = 1'b0;
    assign row1_vec[9] = 1'b0;
    assign row1_vec[10] = 1'b0;
    assign row1_vec[11] = 1'b0;
    assign row1_vec[12] = 1'b0;
    assign row1_vec[13] = 1'b0;
    assign row1_vec[14] = 1'b0;
    assign row1_vec[15] = 1'b0;
    assign row1_vec[16] = 1'b0;
    assign row1_vec[17] = 1'b0;
    assign row1_vec[18] = 1'b0;
    assign row1_vec[19] = 1'b0;
    assign row1_vec[20] = 1'b0;
    assign row1_vec[21] = 1'b0;
    assign row1_vec[22] = 1'b0;
    assign row1_vec[23] = 1'b0;
    assign row1_vec[24] = 1'b0;
    assign row1_vec[25] = 1'b0;
    assign row1_vec[26] = 1'b0;
    assign row1_vec[51] = 1'b0;

    assign p = row0_vec + row1_vec;
endmodule
