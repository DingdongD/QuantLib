
// `include "csa.v"
module wallace_tree_26x24 (
    input [25:0] a,
    input [23:0] b,
    output [49:8] x,  // sum high
    output [49:8] y,  // carry high
    output [7:0] z         // sum low
);

reg [23:0] p [0:25];  // partial products
parameter zero = 1'b0;
integer i,j;
always @* begin
    for(i=0;i<26;i=i+1)
        for(j=0;j<24;j=j+1)
            p[i][j] = a[i] & b[j];
end

wire c_overflow;  // highest carry


// level 0
wire [7:0] s0[0:49];
wire [7:0] c0[0:49];
csa a0_1_0 (p[0][1],p[1][0],zero,s0[1][0],c0[2][0]);
csa a0_2_0 (p[0][2],p[1][1],p[2][0],s0[2][0],c0[3][0]);
csa a0_3_0 (p[0][3],p[1][2],p[2][1],s0[3][0],c0[4][0]);
csa a0_4_0 (p[0][4],p[1][3],p[2][2],s0[4][0],c0[5][0]);
csa a0_4_1 (p[3][1],p[4][0],zero,s0[4][1],c0[5][1]);
csa a0_5_0 (p[0][5],p[1][4],p[2][3],s0[5][0],c0[6][0]);
csa a0_5_1 (p[3][2],p[4][1],p[5][0],s0[5][1],c0[6][1]);
csa a0_6_0 (p[0][6],p[1][5],p[2][4],s0[6][0],c0[7][0]);
csa a0_6_1 (p[3][3],p[4][2],p[5][1],s0[6][1],c0[7][1]);
csa a0_7_0 (p[0][7],p[1][6],p[2][5],s0[7][0],c0[8][0]);
csa a0_7_1 (p[3][4],p[4][3],p[5][2],s0[7][1],c0[8][1]);
csa a0_7_2 (p[6][1],p[7][0],zero,s0[7][2],c0[8][2]);
csa a0_8_0 (p[0][8],p[1][7],p[2][6],s0[8][0],c0[9][0]);
csa a0_8_1 (p[3][5],p[4][4],p[5][3],s0[8][1],c0[9][1]);
csa a0_8_2 (p[6][2],p[7][1],p[8][0],s0[8][2],c0[9][2]);
csa a0_9_0 (p[0][9],p[1][8],p[2][7],s0[9][0],c0[10][0]);
csa a0_9_1 (p[3][6],p[4][5],p[5][4],s0[9][1],c0[10][1]);
csa a0_9_2 (p[6][3],p[7][2],p[8][1],s0[9][2],c0[10][2]);
csa a0_10_0 (p[0][10],p[1][9],p[2][8],s0[10][0],c0[11][0]);
csa a0_10_1 (p[3][7],p[4][6],p[5][5],s0[10][1],c0[11][1]);
csa a0_10_2 (p[6][4],p[7][3],p[8][2],s0[10][2],c0[11][2]);
csa a0_10_3 (p[9][1],p[10][0],zero,s0[10][3],c0[11][3]);
csa a0_11_0 (p[0][11],p[1][10],p[2][9],s0[11][0],c0[12][0]);
csa a0_11_1 (p[3][8],p[4][7],p[5][6],s0[11][1],c0[12][1]);
csa a0_11_2 (p[6][5],p[7][4],p[8][3],s0[11][2],c0[12][2]);
csa a0_11_3 (p[9][2],p[10][1],p[11][0],s0[11][3],c0[12][3]);
csa a0_12_0 (p[0][12],p[1][11],p[2][10],s0[12][0],c0[13][0]);
csa a0_12_1 (p[3][9],p[4][8],p[5][7],s0[12][1],c0[13][1]);
csa a0_12_2 (p[6][6],p[7][5],p[8][4],s0[12][2],c0[13][2]);
csa a0_12_3 (p[9][3],p[10][2],p[11][1],s0[12][3],c0[13][3]);
csa a0_13_0 (p[0][13],p[1][12],p[2][11],s0[13][0],c0[14][0]);
csa a0_13_1 (p[3][10],p[4][9],p[5][8],s0[13][1],c0[14][1]);
csa a0_13_2 (p[6][7],p[7][6],p[8][5],s0[13][2],c0[14][2]);
csa a0_13_3 (p[9][4],p[10][3],p[11][2],s0[13][3],c0[14][3]);
csa a0_13_4 (p[12][1],p[13][0],zero,s0[13][4],c0[14][4]);
csa a0_14_0 (p[0][14],p[1][13],p[2][12],s0[14][0],c0[15][0]);
csa a0_14_1 (p[3][11],p[4][10],p[5][9],s0[14][1],c0[15][1]);
csa a0_14_2 (p[6][8],p[7][7],p[8][6],s0[14][2],c0[15][2]);
csa a0_14_3 (p[9][5],p[10][4],p[11][3],s0[14][3],c0[15][3]);
csa a0_14_4 (p[12][2],p[13][1],p[14][0],s0[14][4],c0[15][4]);
csa a0_15_0 (p[0][15],p[1][14],p[2][13],s0[15][0],c0[16][0]);
csa a0_15_1 (p[3][12],p[4][11],p[5][10],s0[15][1],c0[16][1]);
csa a0_15_2 (p[6][9],p[7][8],p[8][7],s0[15][2],c0[16][2]);
csa a0_15_3 (p[9][6],p[10][5],p[11][4],s0[15][3],c0[16][3]);
csa a0_15_4 (p[12][3],p[13][2],p[14][1],s0[15][4],c0[16][4]);
csa a0_16_0 (p[0][16],p[1][15],p[2][14],s0[16][0],c0[17][0]);
csa a0_16_1 (p[3][13],p[4][12],p[5][11],s0[16][1],c0[17][1]);
csa a0_16_2 (p[6][10],p[7][9],p[8][8],s0[16][2],c0[17][2]);
csa a0_16_3 (p[9][7],p[10][6],p[11][5],s0[16][3],c0[17][3]);
csa a0_16_4 (p[12][4],p[13][3],p[14][2],s0[16][4],c0[17][4]);
csa a0_16_5 (p[15][1],p[16][0],zero,s0[16][5],c0[17][5]);
csa a0_17_0 (p[0][17],p[1][16],p[2][15],s0[17][0],c0[18][0]);
csa a0_17_1 (p[3][14],p[4][13],p[5][12],s0[17][1],c0[18][1]);
csa a0_17_2 (p[6][11],p[7][10],p[8][9],s0[17][2],c0[18][2]);
csa a0_17_3 (p[9][8],p[10][7],p[11][6],s0[17][3],c0[18][3]);
csa a0_17_4 (p[12][5],p[13][4],p[14][3],s0[17][4],c0[18][4]);
csa a0_17_5 (p[15][2],p[16][1],p[17][0],s0[17][5],c0[18][5]);
csa a0_18_0 (p[0][18],p[1][17],p[2][16],s0[18][0],c0[19][0]);
csa a0_18_1 (p[3][15],p[4][14],p[5][13],s0[18][1],c0[19][1]);
csa a0_18_2 (p[6][12],p[7][11],p[8][10],s0[18][2],c0[19][2]);
csa a0_18_3 (p[9][9],p[10][8],p[11][7],s0[18][3],c0[19][3]);
csa a0_18_4 (p[12][6],p[13][5],p[14][4],s0[18][4],c0[19][4]);
csa a0_18_5 (p[15][3],p[16][2],p[17][1],s0[18][5],c0[19][5]);
csa a0_19_0 (p[0][19],p[1][18],p[2][17],s0[19][0],c0[20][0]);
csa a0_19_1 (p[3][16],p[4][15],p[5][14],s0[19][1],c0[20][1]);
csa a0_19_2 (p[6][13],p[7][12],p[8][11],s0[19][2],c0[20][2]);
csa a0_19_3 (p[9][10],p[10][9],p[11][8],s0[19][3],c0[20][3]);
csa a0_19_4 (p[12][7],p[13][6],p[14][5],s0[19][4],c0[20][4]);
csa a0_19_5 (p[15][4],p[16][3],p[17][2],s0[19][5],c0[20][5]);
csa a0_19_6 (p[18][1],p[19][0],zero,s0[19][6],c0[20][6]);
csa a0_20_0 (p[0][20],p[1][19],p[2][18],s0[20][0],c0[21][0]);
csa a0_20_1 (p[3][17],p[4][16],p[5][15],s0[20][1],c0[21][1]);
csa a0_20_2 (p[6][14],p[7][13],p[8][12],s0[20][2],c0[21][2]);
csa a0_20_3 (p[9][11],p[10][10],p[11][9],s0[20][3],c0[21][3]);
csa a0_20_4 (p[12][8],p[13][7],p[14][6],s0[20][4],c0[21][4]);
csa a0_20_5 (p[15][5],p[16][4],p[17][3],s0[20][5],c0[21][5]);
csa a0_20_6 (p[18][2],p[19][1],p[20][0],s0[20][6],c0[21][6]);
csa a0_21_0 (p[0][21],p[1][20],p[2][19],s0[21][0],c0[22][0]);
csa a0_21_1 (p[3][18],p[4][17],p[5][16],s0[21][1],c0[22][1]);
csa a0_21_2 (p[6][15],p[7][14],p[8][13],s0[21][2],c0[22][2]);
csa a0_21_3 (p[9][12],p[10][11],p[11][10],s0[21][3],c0[22][3]);
csa a0_21_4 (p[12][9],p[13][8],p[14][7],s0[21][4],c0[22][4]);
csa a0_21_5 (p[15][6],p[16][5],p[17][4],s0[21][5],c0[22][5]);
csa a0_21_6 (p[18][3],p[19][2],p[20][1],s0[21][6],c0[22][6]);
csa a0_22_0 (p[0][22],p[1][21],p[2][20],s0[22][0],c0[23][0]);
csa a0_22_1 (p[3][19],p[4][18],p[5][17],s0[22][1],c0[23][1]);
csa a0_22_2 (p[6][16],p[7][15],p[8][14],s0[22][2],c0[23][2]);
csa a0_22_3 (p[9][13],p[10][12],p[11][11],s0[22][3],c0[23][3]);
csa a0_22_4 (p[12][10],p[13][9],p[14][8],s0[22][4],c0[23][4]);
csa a0_22_5 (p[15][7],p[16][6],p[17][5],s0[22][5],c0[23][5]);
csa a0_22_6 (p[18][4],p[19][3],p[20][2],s0[22][6],c0[23][6]);
csa a0_22_7 (p[21][1],p[22][0],zero,s0[22][7],c0[23][7]);
csa a0_23_0 (p[0][23],p[1][22],p[2][21],s0[23][0],c0[24][0]);
csa a0_23_1 (p[3][20],p[4][19],p[5][18],s0[23][1],c0[24][1]);
csa a0_23_2 (p[6][17],p[7][16],p[8][15],s0[23][2],c0[24][2]);
csa a0_23_3 (p[9][14],p[10][13],p[11][12],s0[23][3],c0[24][3]);
csa a0_23_4 (p[12][11],p[13][10],p[14][9],s0[23][4],c0[24][4]);
csa a0_23_5 (p[15][8],p[16][7],p[17][6],s0[23][5],c0[24][5]);
csa a0_23_6 (p[18][5],p[19][4],p[20][3],s0[23][6],c0[24][6]);
csa a0_23_7 (p[21][2],p[22][1],p[23][0],s0[23][7],c0[24][7]);
csa a0_24_0 (p[1][23],p[2][22],p[3][21],s0[24][0],c0[25][0]);
csa a0_24_1 (p[4][20],p[5][19],p[6][18],s0[24][1],c0[25][1]);
csa a0_24_2 (p[7][17],p[8][16],p[9][15],s0[24][2],c0[25][2]);
csa a0_24_3 (p[10][14],p[11][13],p[12][12],s0[24][3],c0[25][3]);
csa a0_24_4 (p[13][11],p[14][10],p[15][9],s0[24][4],c0[25][4]);
csa a0_24_5 (p[16][8],p[17][7],p[18][6],s0[24][5],c0[25][5]);
csa a0_24_6 (p[19][5],p[20][4],p[21][3],s0[24][6],c0[25][6]);
csa a0_24_7 (p[22][2],p[23][1],p[24][0],s0[24][7],c0[25][7]);
csa a0_25_0 (p[2][23],p[3][22],p[4][21],s0[25][0],c0[26][0]);
csa a0_25_1 (p[5][20],p[6][19],p[7][18],s0[25][1],c0[26][1]);
csa a0_25_2 (p[8][17],p[9][16],p[10][15],s0[25][2],c0[26][2]);
csa a0_25_3 (p[11][14],p[12][13],p[13][12],s0[25][3],c0[26][3]);
csa a0_25_4 (p[14][11],p[15][10],p[16][9],s0[25][4],c0[26][4]);
csa a0_25_5 (p[17][8],p[18][7],p[19][6],s0[25][5],c0[26][5]);
csa a0_25_6 (p[20][5],p[21][4],p[22][3],s0[25][6],c0[26][6]);
csa a0_25_7 (p[23][2],p[24][1],p[25][0],s0[25][7],c0[26][7]);
csa a0_26_0 (p[3][23],p[4][22],p[5][21],s0[26][0],c0[27][0]);
csa a0_26_1 (p[6][20],p[7][19],p[8][18],s0[26][1],c0[27][1]);
csa a0_26_2 (p[9][17],p[10][16],p[11][15],s0[26][2],c0[27][2]);
csa a0_26_3 (p[12][14],p[13][13],p[14][12],s0[26][3],c0[27][3]);
csa a0_26_4 (p[15][11],p[16][10],p[17][9],s0[26][4],c0[27][4]);
csa a0_26_5 (p[18][8],p[19][7],p[20][6],s0[26][5],c0[27][5]);
csa a0_26_6 (p[21][5],p[22][4],p[23][3],s0[26][6],c0[27][6]);
csa a0_26_7 (p[24][2],p[25][1],zero,s0[26][7],c0[27][7]);
csa a0_27_0 (p[4][23],p[5][22],p[6][21],s0[27][0],c0[28][0]);
csa a0_27_1 (p[7][20],p[8][19],p[9][18],s0[27][1],c0[28][1]);
csa a0_27_2 (p[10][17],p[11][16],p[12][15],s0[27][2],c0[28][2]);
csa a0_27_3 (p[13][14],p[14][13],p[15][12],s0[27][3],c0[28][3]);
csa a0_27_4 (p[16][11],p[17][10],p[18][9],s0[27][4],c0[28][4]);
csa a0_27_5 (p[19][8],p[20][7],p[21][6],s0[27][5],c0[28][5]);
csa a0_27_6 (p[22][5],p[23][4],p[24][3],s0[27][6],c0[28][6]);
csa a0_28_0 (p[5][23],p[6][22],p[7][21],s0[28][0],c0[29][0]);
csa a0_28_1 (p[8][20],p[9][19],p[10][18],s0[28][1],c0[29][1]);
csa a0_28_2 (p[11][17],p[12][16],p[13][15],s0[28][2],c0[29][2]);
csa a0_28_3 (p[14][14],p[15][13],p[16][12],s0[28][3],c0[29][3]);
csa a0_28_4 (p[17][11],p[18][10],p[19][9],s0[28][4],c0[29][4]);
csa a0_28_5 (p[20][8],p[21][7],p[22][6],s0[28][5],c0[29][5]);
csa a0_28_6 (p[23][5],p[24][4],p[25][3],s0[28][6],c0[29][6]);
csa a0_29_0 (p[6][23],p[7][22],p[8][21],s0[29][0],c0[30][0]);
csa a0_29_1 (p[9][20],p[10][19],p[11][18],s0[29][1],c0[30][1]);
csa a0_29_2 (p[12][17],p[13][16],p[14][15],s0[29][2],c0[30][2]);
csa a0_29_3 (p[15][14],p[16][13],p[17][12],s0[29][3],c0[30][3]);
csa a0_29_4 (p[18][11],p[19][10],p[20][9],s0[29][4],c0[30][4]);
csa a0_29_5 (p[21][8],p[22][7],p[23][6],s0[29][5],c0[30][5]);
csa a0_29_6 (p[24][5],p[25][4],zero,s0[29][6],c0[30][6]);
csa a0_30_0 (p[7][23],p[8][22],p[9][21],s0[30][0],c0[31][0]);
csa a0_30_1 (p[10][20],p[11][19],p[12][18],s0[30][1],c0[31][1]);
csa a0_30_2 (p[13][17],p[14][16],p[15][15],s0[30][2],c0[31][2]);
csa a0_30_3 (p[16][14],p[17][13],p[18][12],s0[30][3],c0[31][3]);
csa a0_30_4 (p[19][11],p[20][10],p[21][9],s0[30][4],c0[31][4]);
csa a0_30_5 (p[22][8],p[23][7],p[24][6],s0[30][5],c0[31][5]);
csa a0_31_0 (p[8][23],p[9][22],p[10][21],s0[31][0],c0[32][0]);
csa a0_31_1 (p[11][20],p[12][19],p[13][18],s0[31][1],c0[32][1]);
csa a0_31_2 (p[14][17],p[15][16],p[16][15],s0[31][2],c0[32][2]);
csa a0_31_3 (p[17][14],p[18][13],p[19][12],s0[31][3],c0[32][3]);
csa a0_31_4 (p[20][11],p[21][10],p[22][9],s0[31][4],c0[32][4]);
csa a0_31_5 (p[23][8],p[24][7],p[25][6],s0[31][5],c0[32][5]);
csa a0_32_0 (p[9][23],p[10][22],p[11][21],s0[32][0],c0[33][0]);
csa a0_32_1 (p[12][20],p[13][19],p[14][18],s0[32][1],c0[33][1]);
csa a0_32_2 (p[15][17],p[16][16],p[17][15],s0[32][2],c0[33][2]);
csa a0_32_3 (p[18][14],p[19][13],p[20][12],s0[32][3],c0[33][3]);
csa a0_32_4 (p[21][11],p[22][10],p[23][9],s0[32][4],c0[33][4]);
csa a0_32_5 (p[24][8],p[25][7],zero,s0[32][5],c0[33][5]);
csa a0_33_0 (p[10][23],p[11][22],p[12][21],s0[33][0],c0[34][0]);
csa a0_33_1 (p[13][20],p[14][19],p[15][18],s0[33][1],c0[34][1]);
csa a0_33_2 (p[16][17],p[17][16],p[18][15],s0[33][2],c0[34][2]);
csa a0_33_3 (p[19][14],p[20][13],p[21][12],s0[33][3],c0[34][3]);
csa a0_33_4 (p[22][11],p[23][10],p[24][9],s0[33][4],c0[34][4]);
csa a0_34_0 (p[11][23],p[12][22],p[13][21],s0[34][0],c0[35][0]);
csa a0_34_1 (p[14][20],p[15][19],p[16][18],s0[34][1],c0[35][1]);
csa a0_34_2 (p[17][17],p[18][16],p[19][15],s0[34][2],c0[35][2]);
csa a0_34_3 (p[20][14],p[21][13],p[22][12],s0[34][3],c0[35][3]);
csa a0_34_4 (p[23][11],p[24][10],p[25][9],s0[34][4],c0[35][4]);
csa a0_35_0 (p[12][23],p[13][22],p[14][21],s0[35][0],c0[36][0]);
csa a0_35_1 (p[15][20],p[16][19],p[17][18],s0[35][1],c0[36][1]);
csa a0_35_2 (p[18][17],p[19][16],p[20][15],s0[35][2],c0[36][2]);
csa a0_35_3 (p[21][14],p[22][13],p[23][12],s0[35][3],c0[36][3]);
csa a0_35_4 (p[24][11],p[25][10],zero,s0[35][4],c0[36][4]);
csa a0_36_0 (p[13][23],p[14][22],p[15][21],s0[36][0],c0[37][0]);
csa a0_36_1 (p[16][20],p[17][19],p[18][18],s0[36][1],c0[37][1]);
csa a0_36_2 (p[19][17],p[20][16],p[21][15],s0[36][2],c0[37][2]);
csa a0_36_3 (p[22][14],p[23][13],p[24][12],s0[36][3],c0[37][3]);
csa a0_37_0 (p[14][23],p[15][22],p[16][21],s0[37][0],c0[38][0]);
csa a0_37_1 (p[17][20],p[18][19],p[19][18],s0[37][1],c0[38][1]);
csa a0_37_2 (p[20][17],p[21][16],p[22][15],s0[37][2],c0[38][2]);
csa a0_37_3 (p[23][14],p[24][13],p[25][12],s0[37][3],c0[38][3]);
csa a0_38_0 (p[15][23],p[16][22],p[17][21],s0[38][0],c0[39][0]);
csa a0_38_1 (p[18][20],p[19][19],p[20][18],s0[38][1],c0[39][1]);
csa a0_38_2 (p[21][17],p[22][16],p[23][15],s0[38][2],c0[39][2]);
csa a0_38_3 (p[24][14],p[25][13],zero,s0[38][3],c0[39][3]);
csa a0_39_0 (p[16][23],p[17][22],p[18][21],s0[39][0],c0[40][0]);
csa a0_39_1 (p[19][20],p[20][19],p[21][18],s0[39][1],c0[40][1]);
csa a0_39_2 (p[22][17],p[23][16],p[24][15],s0[39][2],c0[40][2]);
csa a0_40_0 (p[17][23],p[18][22],p[19][21],s0[40][0],c0[41][0]);
csa a0_40_1 (p[20][20],p[21][19],p[22][18],s0[40][1],c0[41][1]);
csa a0_40_2 (p[23][17],p[24][16],p[25][15],s0[40][2],c0[41][2]);
csa a0_41_0 (p[18][23],p[19][22],p[20][21],s0[41][0],c0[42][0]);
csa a0_41_1 (p[21][20],p[22][19],p[23][18],s0[41][1],c0[42][1]);
csa a0_41_2 (p[24][17],p[25][16],zero,s0[41][2],c0[42][2]);
csa a0_42_0 (p[19][23],p[20][22],p[21][21],s0[42][0],c0[43][0]);
csa a0_42_1 (p[22][20],p[23][19],p[24][18],s0[42][1],c0[43][1]);
csa a0_43_0 (p[20][23],p[21][22],p[22][21],s0[43][0],c0[44][0]);
csa a0_43_1 (p[23][20],p[24][19],p[25][18],s0[43][1],c0[44][1]);
csa a0_44_0 (p[21][23],p[22][22],p[23][21],s0[44][0],c0[45][0]);
csa a0_44_1 (p[24][20],p[25][19],zero,s0[44][1],c0[45][1]);
csa a0_45_0 (p[22][23],p[23][22],p[24][21],s0[45][0],c0[46][0]);
csa a0_46_0 (p[23][23],p[24][22],p[25][21],s0[46][0],c0[47][0]);
csa a0_47_0 (p[24][23],p[25][22],zero,s0[47][0],c0[48][0]);

// level 1
wire [4:0] s1[0:49];
wire [4:0] c1[0:49];
csa a1_2_0 (c0[2][0],s0[2][0],zero,s1[2][0],c1[3][0]);
csa a1_3_0 (c0[3][0],s0[3][0],p[3][0],s1[3][0],c1[4][0]);
csa a1_4_0 (c0[4][0],s0[4][0],s0[4][1],s1[4][0],c1[5][0]);
csa a1_5_0 (c0[5][0],c0[5][1],s0[5][0],s1[5][0],c1[6][0]);
csa a1_6_0 (c0[6][0],c0[6][1],s0[6][0],s1[6][0],c1[7][0]);
csa a1_6_1 (s0[6][1],p[6][0],zero,s1[6][1],c1[7][1]);
csa a1_7_0 (c0[7][0],c0[7][1],s0[7][0],s1[7][0],c1[8][0]);
csa a1_7_1 (s0[7][1],s0[7][2],zero,s1[7][1],c1[8][1]);
csa a1_8_0 (c0[8][0],c0[8][1],c0[8][2],s1[8][0],c1[9][0]);
csa a1_8_1 (s0[8][0],s0[8][1],s0[8][2],s1[8][1],c1[9][1]);
csa a1_9_0 (c0[9][0],c0[9][1],c0[9][2],s1[9][0],c1[10][0]);
csa a1_9_1 (s0[9][0],s0[9][1],s0[9][2],s1[9][1],c1[10][1]);
csa a1_10_0 (c0[10][0],c0[10][1],c0[10][2],s1[10][0],c1[11][0]);
csa a1_10_1 (s0[10][0],s0[10][1],s0[10][2],s1[10][1],c1[11][1]);
csa a1_11_0 (c0[11][0],c0[11][1],c0[11][2],s1[11][0],c1[12][0]);
csa a1_11_1 (c0[11][3],s0[11][0],s0[11][1],s1[11][1],c1[12][1]);
csa a1_11_2 (s0[11][2],s0[11][3],zero,s1[11][2],c1[12][2]);
csa a1_12_0 (c0[12][0],c0[12][1],c0[12][2],s1[12][0],c1[13][0]);
csa a1_12_1 (c0[12][3],s0[12][0],s0[12][1],s1[12][1],c1[13][1]);
csa a1_12_2 (s0[12][2],s0[12][3],p[12][0],s1[12][2],c1[13][2]);
csa a1_13_0 (c0[13][0],c0[13][1],c0[13][2],s1[13][0],c1[14][0]);
csa a1_13_1 (c0[13][3],s0[13][0],s0[13][1],s1[13][1],c1[14][1]);
csa a1_13_2 (s0[13][2],s0[13][3],s0[13][4],s1[13][2],c1[14][2]);
csa a1_14_0 (c0[14][0],c0[14][1],c0[14][2],s1[14][0],c1[15][0]);
csa a1_14_1 (c0[14][3],c0[14][4],s0[14][0],s1[14][1],c1[15][1]);
csa a1_14_2 (s0[14][1],s0[14][2],s0[14][3],s1[14][2],c1[15][2]);
csa a1_15_0 (c0[15][0],c0[15][1],c0[15][2],s1[15][0],c1[16][0]);
csa a1_15_1 (c0[15][3],c0[15][4],s0[15][0],s1[15][1],c1[16][1]);
csa a1_15_2 (s0[15][1],s0[15][2],s0[15][3],s1[15][2],c1[16][2]);
csa a1_15_3 (s0[15][4],p[15][0],zero,s1[15][3],c1[16][3]);
csa a1_16_0 (c0[16][0],c0[16][1],c0[16][2],s1[16][0],c1[17][0]);
csa a1_16_1 (c0[16][3],c0[16][4],s0[16][0],s1[16][1],c1[17][1]);
csa a1_16_2 (s0[16][1],s0[16][2],s0[16][3],s1[16][2],c1[17][2]);
csa a1_16_3 (s0[16][4],s0[16][5],zero,s1[16][3],c1[17][3]);
csa a1_17_0 (c0[17][0],c0[17][1],c0[17][2],s1[17][0],c1[18][0]);
csa a1_17_1 (c0[17][3],c0[17][4],c0[17][5],s1[17][1],c1[18][1]);
csa a1_17_2 (s0[17][0],s0[17][1],s0[17][2],s1[17][2],c1[18][2]);
csa a1_17_3 (s0[17][3],s0[17][4],s0[17][5],s1[17][3],c1[18][3]);
csa a1_18_0 (c0[18][0],c0[18][1],c0[18][2],s1[18][0],c1[19][0]);
csa a1_18_1 (c0[18][3],c0[18][4],c0[18][5],s1[18][1],c1[19][1]);
csa a1_18_2 (s0[18][0],s0[18][1],s0[18][2],s1[18][2],c1[19][2]);
csa a1_18_3 (s0[18][3],s0[18][4],s0[18][5],s1[18][3],c1[19][3]);
csa a1_19_0 (c0[19][0],c0[19][1],c0[19][2],s1[19][0],c1[20][0]);
csa a1_19_1 (c0[19][3],c0[19][4],c0[19][5],s1[19][1],c1[20][1]);
csa a1_19_2 (s0[19][0],s0[19][1],s0[19][2],s1[19][2],c1[20][2]);
csa a1_19_3 (s0[19][3],s0[19][4],s0[19][5],s1[19][3],c1[20][3]);
csa a1_20_0 (c0[20][0],c0[20][1],c0[20][2],s1[20][0],c1[21][0]);
csa a1_20_1 (c0[20][3],c0[20][4],c0[20][5],s1[20][1],c1[21][1]);
csa a1_20_2 (c0[20][6],s0[20][0],s0[20][1],s1[20][2],c1[21][2]);
csa a1_20_3 (s0[20][2],s0[20][3],s0[20][4],s1[20][3],c1[21][3]);
csa a1_20_4 (s0[20][5],s0[20][6],zero,s1[20][4],c1[21][4]);
csa a1_21_0 (c0[21][0],c0[21][1],c0[21][2],s1[21][0],c1[22][0]);
csa a1_21_1 (c0[21][3],c0[21][4],c0[21][5],s1[21][1],c1[22][1]);
csa a1_21_2 (c0[21][6],s0[21][0],s0[21][1],s1[21][2],c1[22][2]);
csa a1_21_3 (s0[21][2],s0[21][3],s0[21][4],s1[21][3],c1[22][3]);
csa a1_21_4 (s0[21][5],s0[21][6],p[21][0],s1[21][4],c1[22][4]);
csa a1_22_0 (c0[22][0],c0[22][1],c0[22][2],s1[22][0],c1[23][0]);
csa a1_22_1 (c0[22][3],c0[22][4],c0[22][5],s1[22][1],c1[23][1]);
csa a1_22_2 (c0[22][6],s0[22][0],s0[22][1],s1[22][2],c1[23][2]);
csa a1_22_3 (s0[22][2],s0[22][3],s0[22][4],s1[22][3],c1[23][3]);
csa a1_22_4 (s0[22][5],s0[22][6],s0[22][7],s1[22][4],c1[23][4]);
csa a1_23_0 (c0[23][0],c0[23][1],c0[23][2],s1[23][0],c1[24][0]);
csa a1_23_1 (c0[23][3],c0[23][4],c0[23][5],s1[23][1],c1[24][1]);
csa a1_23_2 (c0[23][6],c0[23][7],s0[23][0],s1[23][2],c1[24][2]);
csa a1_23_3 (s0[23][1],s0[23][2],s0[23][3],s1[23][3],c1[24][3]);
csa a1_23_4 (s0[23][4],s0[23][5],s0[23][6],s1[23][4],c1[24][4]);
csa a1_24_0 (c0[24][0],c0[24][1],c0[24][2],s1[24][0],c1[25][0]);
csa a1_24_1 (c0[24][3],c0[24][4],c0[24][5],s1[24][1],c1[25][1]);
csa a1_24_2 (c0[24][6],c0[24][7],s0[24][0],s1[24][2],c1[25][2]);
csa a1_24_3 (s0[24][1],s0[24][2],s0[24][3],s1[24][3],c1[25][3]);
csa a1_24_4 (s0[24][4],s0[24][5],s0[24][6],s1[24][4],c1[25][4]);
csa a1_25_0 (c0[25][0],c0[25][1],c0[25][2],s1[25][0],c1[26][0]);
csa a1_25_1 (c0[25][3],c0[25][4],c0[25][5],s1[25][1],c1[26][1]);
csa a1_25_2 (c0[25][6],c0[25][7],s0[25][0],s1[25][2],c1[26][2]);
csa a1_25_3 (s0[25][1],s0[25][2],s0[25][3],s1[25][3],c1[26][3]);
csa a1_25_4 (s0[25][4],s0[25][5],s0[25][6],s1[25][4],c1[26][4]);
csa a1_26_0 (c0[26][0],c0[26][1],c0[26][2],s1[26][0],c1[27][0]);
csa a1_26_1 (c0[26][3],c0[26][4],c0[26][5],s1[26][1],c1[27][1]);
csa a1_26_2 (c0[26][6],c0[26][7],s0[26][0],s1[26][2],c1[27][2]);
csa a1_26_3 (s0[26][1],s0[26][2],s0[26][3],s1[26][3],c1[27][3]);
csa a1_26_4 (s0[26][4],s0[26][5],s0[26][6],s1[26][4],c1[27][4]);
csa a1_27_0 (c0[27][0],c0[27][1],c0[27][2],s1[27][0],c1[28][0]);
csa a1_27_1 (c0[27][3],c0[27][4],c0[27][5],s1[27][1],c1[28][1]);
csa a1_27_2 (c0[27][6],c0[27][7],s0[27][0],s1[27][2],c1[28][2]);
csa a1_27_3 (s0[27][1],s0[27][2],s0[27][3],s1[27][3],c1[28][3]);
csa a1_27_4 (s0[27][4],s0[27][5],s0[27][6],s1[27][4],c1[28][4]);
csa a1_28_0 (c0[28][0],c0[28][1],c0[28][2],s1[28][0],c1[29][0]);
csa a1_28_1 (c0[28][3],c0[28][4],c0[28][5],s1[28][1],c1[29][1]);
csa a1_28_2 (c0[28][6],s0[28][0],s0[28][1],s1[28][2],c1[29][2]);
csa a1_28_3 (s0[28][2],s0[28][3],s0[28][4],s1[28][3],c1[29][3]);
csa a1_28_4 (s0[28][5],s0[28][6],zero,s1[28][4],c1[29][4]);
csa a1_29_0 (c0[29][0],c0[29][1],c0[29][2],s1[29][0],c1[30][0]);
csa a1_29_1 (c0[29][3],c0[29][4],c0[29][5],s1[29][1],c1[30][1]);
csa a1_29_2 (c0[29][6],s0[29][0],s0[29][1],s1[29][2],c1[30][2]);
csa a1_29_3 (s0[29][2],s0[29][3],s0[29][4],s1[29][3],c1[30][3]);
csa a1_29_4 (s0[29][5],s0[29][6],zero,s1[29][4],c1[30][4]);
csa a1_30_0 (c0[30][0],c0[30][1],c0[30][2],s1[30][0],c1[31][0]);
csa a1_30_1 (c0[30][3],c0[30][4],c0[30][5],s1[30][1],c1[31][1]);
csa a1_30_2 (c0[30][6],s0[30][0],s0[30][1],s1[30][2],c1[31][2]);
csa a1_30_3 (s0[30][2],s0[30][3],s0[30][4],s1[30][3],c1[31][3]);
csa a1_30_4 (s0[30][5],p[25][5],zero,s1[30][4],c1[31][4]);
csa a1_31_0 (c0[31][0],c0[31][1],c0[31][2],s1[31][0],c1[32][0]);
csa a1_31_1 (c0[31][3],c0[31][4],c0[31][5],s1[31][1],c1[32][1]);
csa a1_31_2 (s0[31][0],s0[31][1],s0[31][2],s1[31][2],c1[32][2]);
csa a1_31_3 (s0[31][3],s0[31][4],s0[31][5],s1[31][3],c1[32][3]);
csa a1_32_0 (c0[32][0],c0[32][1],c0[32][2],s1[32][0],c1[33][0]);
csa a1_32_1 (c0[32][3],c0[32][4],c0[32][5],s1[32][1],c1[33][1]);
csa a1_32_2 (s0[32][0],s0[32][1],s0[32][2],s1[32][2],c1[33][2]);
csa a1_32_3 (s0[32][3],s0[32][4],s0[32][5],s1[32][3],c1[33][3]);
csa a1_33_0 (c0[33][0],c0[33][1],c0[33][2],s1[33][0],c1[34][0]);
csa a1_33_1 (c0[33][3],c0[33][4],c0[33][5],s1[33][1],c1[34][1]);
csa a1_33_2 (s0[33][0],s0[33][1],s0[33][2],s1[33][2],c1[34][2]);
csa a1_33_3 (s0[33][3],s0[33][4],p[25][8],s1[33][3],c1[34][3]);
csa a1_34_0 (c0[34][0],c0[34][1],c0[34][2],s1[34][0],c1[35][0]);
csa a1_34_1 (c0[34][3],c0[34][4],s0[34][0],s1[34][1],c1[35][1]);
csa a1_34_2 (s0[34][1],s0[34][2],s0[34][3],s1[34][2],c1[35][2]);
csa a1_35_0 (c0[35][0],c0[35][1],c0[35][2],s1[35][0],c1[36][0]);
csa a1_35_1 (c0[35][3],c0[35][4],s0[35][0],s1[35][1],c1[36][1]);
csa a1_35_2 (s0[35][1],s0[35][2],s0[35][3],s1[35][2],c1[36][2]);
csa a1_36_0 (c0[36][0],c0[36][1],c0[36][2],s1[36][0],c1[37][0]);
csa a1_36_1 (c0[36][3],c0[36][4],s0[36][0],s1[36][1],c1[37][1]);
csa a1_36_2 (s0[36][1],s0[36][2],s0[36][3],s1[36][2],c1[37][2]);
csa a1_37_0 (c0[37][0],c0[37][1],c0[37][2],s1[37][0],c1[38][0]);
csa a1_37_1 (c0[37][3],s0[37][0],s0[37][1],s1[37][1],c1[38][1]);
csa a1_37_2 (s0[37][2],s0[37][3],zero,s1[37][2],c1[38][2]);
csa a1_38_0 (c0[38][0],c0[38][1],c0[38][2],s1[38][0],c1[39][0]);
csa a1_38_1 (c0[38][3],s0[38][0],s0[38][1],s1[38][1],c1[39][1]);
csa a1_38_2 (s0[38][2],s0[38][3],zero,s1[38][2],c1[39][2]);
csa a1_39_0 (c0[39][0],c0[39][1],c0[39][2],s1[39][0],c1[40][0]);
csa a1_39_1 (c0[39][3],s0[39][0],s0[39][1],s1[39][1],c1[40][1]);
csa a1_39_2 (s0[39][2],p[25][14],zero,s1[39][2],c1[40][2]);
csa a1_40_0 (c0[40][0],c0[40][1],c0[40][2],s1[40][0],c1[41][0]);
csa a1_40_1 (s0[40][0],s0[40][1],s0[40][2],s1[40][1],c1[41][1]);
csa a1_41_0 (c0[41][0],c0[41][1],c0[41][2],s1[41][0],c1[42][0]);
csa a1_41_1 (s0[41][0],s0[41][1],s0[41][2],s1[41][1],c1[42][1]);
csa a1_42_0 (c0[42][0],c0[42][1],c0[42][2],s1[42][0],c1[43][0]);
csa a1_42_1 (s0[42][0],s0[42][1],p[25][17],s1[42][1],c1[43][1]);
csa a1_43_0 (c0[43][0],c0[43][1],s0[43][0],s1[43][0],c1[44][0]);
csa a1_44_0 (c0[44][0],c0[44][1],s0[44][0],s1[44][0],c1[45][0]);
csa a1_45_0 (c0[45][0],c0[45][1],s0[45][0],s1[45][0],c1[46][0]);
csa a1_46_0 (c0[46][0],s0[46][0],zero,s1[46][0],c1[47][0]);
csa a1_47_0 (c0[47][0],s0[47][0],zero,s1[47][0],c1[48][0]);
csa a1_48_0 (c0[48][0],p[25][23],zero,s1[48][0],c1[49][0]);

// level 2
wire [3:0] s2[0:49];
wire [3:0] c2[0:49];
csa a2_3_0 (c1[3][0],s1[3][0],zero,s2[3][0],c2[4][0]);
csa a2_4_0 (c1[4][0],s1[4][0],zero,s2[4][0],c2[5][0]);
csa a2_5_0 (c1[5][0],s1[5][0],s0[5][1],s2[5][0],c2[6][0]);
csa a2_6_0 (c1[6][0],s1[6][0],s1[6][1],s2[6][0],c2[7][0]);
csa a2_7_0 (c1[7][0],c1[7][1],s1[7][0],s2[7][0],c2[8][0]);
csa a2_8_0 (c1[8][0],c1[8][1],s1[8][0],s2[8][0],c2[9][0]);
csa a2_9_0 (c1[9][0],c1[9][1],s1[9][0],s2[9][0],c2[10][0]);
csa a2_9_1 (s1[9][1],p[9][0],zero,s2[9][1],c2[10][1]);
csa a2_10_0 (c1[10][0],c1[10][1],s1[10][0],s2[10][0],c2[11][0]);
csa a2_10_1 (s1[10][1],s0[10][3],zero,s2[10][1],c2[11][1]);
csa a2_11_0 (c1[11][0],c1[11][1],s1[11][0],s2[11][0],c2[12][0]);
csa a2_11_1 (s1[11][1],s1[11][2],zero,s2[11][1],c2[12][1]);
csa a2_12_0 (c1[12][0],c1[12][1],c1[12][2],s2[12][0],c2[13][0]);
csa a2_12_1 (s1[12][0],s1[12][1],s1[12][2],s2[12][1],c2[13][1]);
csa a2_13_0 (c1[13][0],c1[13][1],c1[13][2],s2[13][0],c2[14][0]);
csa a2_13_1 (s1[13][0],s1[13][1],s1[13][2],s2[13][1],c2[14][1]);
csa a2_14_0 (c1[14][0],c1[14][1],c1[14][2],s2[14][0],c2[15][0]);
csa a2_14_1 (s1[14][0],s1[14][1],s1[14][2],s2[14][1],c2[15][1]);
csa a2_15_0 (c1[15][0],c1[15][1],c1[15][2],s2[15][0],c2[16][0]);
csa a2_15_1 (s1[15][0],s1[15][1],s1[15][2],s2[15][1],c2[16][1]);
csa a2_16_0 (c1[16][0],c1[16][1],c1[16][2],s2[16][0],c2[17][0]);
csa a2_16_1 (c1[16][3],s1[16][0],s1[16][1],s2[16][1],c2[17][1]);
csa a2_16_2 (s1[16][2],s1[16][3],zero,s2[16][2],c2[17][2]);
csa a2_17_0 (c1[17][0],c1[17][1],c1[17][2],s2[17][0],c2[18][0]);
csa a2_17_1 (c1[17][3],s1[17][0],s1[17][1],s2[17][1],c2[18][1]);
csa a2_17_2 (s1[17][2],s1[17][3],zero,s2[17][2],c2[18][2]);
csa a2_18_0 (c1[18][0],c1[18][1],c1[18][2],s2[18][0],c2[19][0]);
csa a2_18_1 (c1[18][3],s1[18][0],s1[18][1],s2[18][1],c2[19][1]);
csa a2_18_2 (s1[18][2],s1[18][3],p[18][0],s2[18][2],c2[19][2]);
csa a2_19_0 (c1[19][0],c1[19][1],c1[19][2],s2[19][0],c2[20][0]);
csa a2_19_1 (c1[19][3],s1[19][0],s1[19][1],s2[19][1],c2[20][1]);
csa a2_19_2 (s1[19][2],s1[19][3],s0[19][6],s2[19][2],c2[20][2]);
csa a2_20_0 (c1[20][0],c1[20][1],c1[20][2],s2[20][0],c2[21][0]);
csa a2_20_1 (c1[20][3],s1[20][0],s1[20][1],s2[20][1],c2[21][1]);
csa a2_20_2 (s1[20][2],s1[20][3],s1[20][4],s2[20][2],c2[21][2]);
csa a2_21_0 (c1[21][0],c1[21][1],c1[21][2],s2[21][0],c2[22][0]);
csa a2_21_1 (c1[21][3],c1[21][4],s1[21][0],s2[21][1],c2[22][1]);
csa a2_21_2 (s1[21][1],s1[21][2],s1[21][3],s2[21][2],c2[22][2]);
csa a2_22_0 (c1[22][0],c1[22][1],c1[22][2],s2[22][0],c2[23][0]);
csa a2_22_1 (c1[22][3],c1[22][4],s1[22][0],s2[22][1],c2[23][1]);
csa a2_22_2 (s1[22][1],s1[22][2],s1[22][3],s2[22][2],c2[23][2]);
csa a2_23_0 (c1[23][0],c1[23][1],c1[23][2],s2[23][0],c2[24][0]);
csa a2_23_1 (c1[23][3],c1[23][4],s1[23][0],s2[23][1],c2[24][1]);
csa a2_23_2 (s1[23][1],s1[23][2],s1[23][3],s2[23][2],c2[24][2]);
csa a2_23_3 (s1[23][4],s0[23][7],zero,s2[23][3],c2[24][3]);
csa a2_24_0 (c1[24][0],c1[24][1],c1[24][2],s2[24][0],c2[25][0]);
csa a2_24_1 (c1[24][3],c1[24][4],s1[24][0],s2[24][1],c2[25][1]);
csa a2_24_2 (s1[24][1],s1[24][2],s1[24][3],s2[24][2],c2[25][2]);
csa a2_24_3 (s1[24][4],s0[24][7],zero,s2[24][3],c2[25][3]);
csa a2_25_0 (c1[25][0],c1[25][1],c1[25][2],s2[25][0],c2[26][0]);
csa a2_25_1 (c1[25][3],c1[25][4],s1[25][0],s2[25][1],c2[26][1]);
csa a2_25_2 (s1[25][1],s1[25][2],s1[25][3],s2[25][2],c2[26][2]);
csa a2_25_3 (s1[25][4],s0[25][7],zero,s2[25][3],c2[26][3]);
csa a2_26_0 (c1[26][0],c1[26][1],c1[26][2],s2[26][0],c2[27][0]);
csa a2_26_1 (c1[26][3],c1[26][4],s1[26][0],s2[26][1],c2[27][1]);
csa a2_26_2 (s1[26][1],s1[26][2],s1[26][3],s2[26][2],c2[27][2]);
csa a2_26_3 (s1[26][4],s0[26][7],zero,s2[26][3],c2[27][3]);
csa a2_27_0 (c1[27][0],c1[27][1],c1[27][2],s2[27][0],c2[28][0]);
csa a2_27_1 (c1[27][3],c1[27][4],s1[27][0],s2[27][1],c2[28][1]);
csa a2_27_2 (s1[27][1],s1[27][2],s1[27][3],s2[27][2],c2[28][2]);
csa a2_27_3 (s1[27][4],p[25][2],zero,s2[27][3],c2[28][3]);
csa a2_28_0 (c1[28][0],c1[28][1],c1[28][2],s2[28][0],c2[29][0]);
csa a2_28_1 (c1[28][3],c1[28][4],s1[28][0],s2[28][1],c2[29][1]);
csa a2_28_2 (s1[28][1],s1[28][2],s1[28][3],s2[28][2],c2[29][2]);
csa a2_29_0 (c1[29][0],c1[29][1],c1[29][2],s2[29][0],c2[30][0]);
csa a2_29_1 (c1[29][3],c1[29][4],s1[29][0],s2[29][1],c2[30][1]);
csa a2_29_2 (s1[29][1],s1[29][2],s1[29][3],s2[29][2],c2[30][2]);
csa a2_30_0 (c1[30][0],c1[30][1],c1[30][2],s2[30][0],c2[31][0]);
csa a2_30_1 (c1[30][3],c1[30][4],s1[30][0],s2[30][1],c2[31][1]);
csa a2_30_2 (s1[30][1],s1[30][2],s1[30][3],s2[30][2],c2[31][2]);
csa a2_31_0 (c1[31][0],c1[31][1],c1[31][2],s2[31][0],c2[32][0]);
csa a2_31_1 (c1[31][3],c1[31][4],s1[31][0],s2[31][1],c2[32][1]);
csa a2_31_2 (s1[31][1],s1[31][2],s1[31][3],s2[31][2],c2[32][2]);
csa a2_32_0 (c1[32][0],c1[32][1],c1[32][2],s2[32][0],c2[33][0]);
csa a2_32_1 (c1[32][3],s1[32][0],s1[32][1],s2[32][1],c2[33][1]);
csa a2_32_2 (s1[32][2],s1[32][3],zero,s2[32][2],c2[33][2]);
csa a2_33_0 (c1[33][0],c1[33][1],c1[33][2],s2[33][0],c2[34][0]);
csa a2_33_1 (c1[33][3],s1[33][0],s1[33][1],s2[33][1],c2[34][1]);
csa a2_33_2 (s1[33][2],s1[33][3],zero,s2[33][2],c2[34][2]);
csa a2_34_0 (c1[34][0],c1[34][1],c1[34][2],s2[34][0],c2[35][0]);
csa a2_34_1 (c1[34][3],s1[34][0],s1[34][1],s2[34][1],c2[35][1]);
csa a2_34_2 (s1[34][2],s0[34][4],zero,s2[34][2],c2[35][2]);
csa a2_35_0 (c1[35][0],c1[35][1],c1[35][2],s2[35][0],c2[36][0]);
csa a2_35_1 (s1[35][0],s1[35][1],s1[35][2],s2[35][1],c2[36][1]);
csa a2_36_0 (c1[36][0],c1[36][1],c1[36][2],s2[36][0],c2[37][0]);
csa a2_36_1 (s1[36][0],s1[36][1],s1[36][2],s2[36][1],c2[37][1]);
csa a2_37_0 (c1[37][0],c1[37][1],c1[37][2],s2[37][0],c2[38][0]);
csa a2_37_1 (s1[37][0],s1[37][1],s1[37][2],s2[37][1],c2[38][1]);
csa a2_38_0 (c1[38][0],c1[38][1],c1[38][2],s2[38][0],c2[39][0]);
csa a2_38_1 (s1[38][0],s1[38][1],s1[38][2],s2[38][1],c2[39][1]);
csa a2_39_0 (c1[39][0],c1[39][1],c1[39][2],s2[39][0],c2[40][0]);
csa a2_39_1 (s1[39][0],s1[39][1],s1[39][2],s2[39][1],c2[40][1]);
csa a2_40_0 (c1[40][0],c1[40][1],c1[40][2],s2[40][0],c2[41][0]);
csa a2_40_1 (s1[40][0],s1[40][1],zero,s2[40][1],c2[41][1]);
csa a2_41_0 (c1[41][0],c1[41][1],s1[41][0],s2[41][0],c2[42][0]);
csa a2_42_0 (c1[42][0],c1[42][1],s1[42][0],s2[42][0],c2[43][0]);
csa a2_43_0 (c1[43][0],c1[43][1],s1[43][0],s2[43][0],c2[44][0]);
csa a2_44_0 (c1[44][0],s1[44][0],s0[44][1],s2[44][0],c2[45][0]);
csa a2_45_0 (c1[45][0],s1[45][0],p[25][20],s2[45][0],c2[46][0]);
csa a2_46_0 (c1[46][0],s1[46][0],zero,s2[46][0],c2[47][0]);
csa a2_47_0 (c1[47][0],s1[47][0],zero,s2[47][0],c2[48][0]);
csa a2_48_0 (c1[48][0],s1[48][0],zero,s2[48][0],c2[49][0]);

// level 3
wire [2:0] s3[0:49];
wire [2:0] c3[0:49];
csa a3_4_0 (c2[4][0],s2[4][0],zero,s3[4][0],c3[5][0]);
csa a3_5_0 (c2[5][0],s2[5][0],zero,s3[5][0],c3[6][0]);
csa a3_6_0 (c2[6][0],s2[6][0],zero,s3[6][0],c3[7][0]);
csa a3_7_0 (c2[7][0],s2[7][0],s1[7][1],s3[7][0],c3[8][0]);
csa a3_8_0 (c2[8][0],s2[8][0],s1[8][1],s3[8][0],c3[9][0]);
csa a3_9_0 (c2[9][0],s2[9][0],s2[9][1],s3[9][0],c3[10][0]);
csa a3_10_0 (c2[10][0],c2[10][1],s2[10][0],s3[10][0],c3[11][0]);
csa a3_11_0 (c2[11][0],c2[11][1],s2[11][0],s3[11][0],c3[12][0]);
csa a3_12_0 (c2[12][0],c2[12][1],s2[12][0],s3[12][0],c3[13][0]);
csa a3_13_0 (c2[13][0],c2[13][1],s2[13][0],s3[13][0],c3[14][0]);
csa a3_14_0 (c2[14][0],c2[14][1],s2[14][0],s3[14][0],c3[15][0]);
csa a3_14_1 (s2[14][1],s0[14][4],zero,s3[14][1],c3[15][1]);
csa a3_15_0 (c2[15][0],c2[15][1],s2[15][0],s3[15][0],c3[16][0]);
csa a3_15_1 (s2[15][1],s1[15][3],zero,s3[15][1],c3[16][1]);
csa a3_16_0 (c2[16][0],c2[16][1],s2[16][0],s3[16][0],c3[17][0]);
csa a3_16_1 (s2[16][1],s2[16][2],zero,s3[16][1],c3[17][1]);
csa a3_17_0 (c2[17][0],c2[17][1],c2[17][2],s3[17][0],c3[18][0]);
csa a3_17_1 (s2[17][0],s2[17][1],s2[17][2],s3[17][1],c3[18][1]);
csa a3_18_0 (c2[18][0],c2[18][1],c2[18][2],s3[18][0],c3[19][0]);
csa a3_18_1 (s2[18][0],s2[18][1],s2[18][2],s3[18][1],c3[19][1]);
csa a3_19_0 (c2[19][0],c2[19][1],c2[19][2],s3[19][0],c3[20][0]);
csa a3_19_1 (s2[19][0],s2[19][1],s2[19][2],s3[19][1],c3[20][1]);
csa a3_20_0 (c2[20][0],c2[20][1],c2[20][2],s3[20][0],c3[21][0]);
csa a3_20_1 (s2[20][0],s2[20][1],s2[20][2],s3[20][1],c3[21][1]);
csa a3_21_0 (c2[21][0],c2[21][1],c2[21][2],s3[21][0],c3[22][0]);
csa a3_21_1 (s2[21][0],s2[21][1],s2[21][2],s3[21][1],c3[22][1]);
csa a3_22_0 (c2[22][0],c2[22][1],c2[22][2],s3[22][0],c3[23][0]);
csa a3_22_1 (s2[22][0],s2[22][1],s2[22][2],s3[22][1],c3[23][1]);
csa a3_23_0 (c2[23][0],c2[23][1],c2[23][2],s3[23][0],c3[24][0]);
csa a3_23_1 (s2[23][0],s2[23][1],s2[23][2],s3[23][1],c3[24][1]);
csa a3_24_0 (c2[24][0],c2[24][1],c2[24][2],s3[24][0],c3[25][0]);
csa a3_24_1 (c2[24][3],s2[24][0],s2[24][1],s3[24][1],c3[25][1]);
csa a3_24_2 (s2[24][2],s2[24][3],zero,s3[24][2],c3[25][2]);
csa a3_25_0 (c2[25][0],c2[25][1],c2[25][2],s3[25][0],c3[26][0]);
csa a3_25_1 (c2[25][3],s2[25][0],s2[25][1],s3[25][1],c3[26][1]);
csa a3_25_2 (s2[25][2],s2[25][3],zero,s3[25][2],c3[26][2]);
csa a3_26_0 (c2[26][0],c2[26][1],c2[26][2],s3[26][0],c3[27][0]);
csa a3_26_1 (c2[26][3],s2[26][0],s2[26][1],s3[26][1],c3[27][1]);
csa a3_26_2 (s2[26][2],s2[26][3],zero,s3[26][2],c3[27][2]);
csa a3_27_0 (c2[27][0],c2[27][1],c2[27][2],s3[27][0],c3[28][0]);
csa a3_27_1 (c2[27][3],s2[27][0],s2[27][1],s3[27][1],c3[28][1]);
csa a3_27_2 (s2[27][2],s2[27][3],zero,s3[27][2],c3[28][2]);
csa a3_28_0 (c2[28][0],c2[28][1],c2[28][2],s3[28][0],c3[29][0]);
csa a3_28_1 (c2[28][3],s2[28][0],s2[28][1],s3[28][1],c3[29][1]);
csa a3_28_2 (s2[28][2],s1[28][4],zero,s3[28][2],c3[29][2]);
csa a3_29_0 (c2[29][0],c2[29][1],c2[29][2],s3[29][0],c3[30][0]);
csa a3_29_1 (s2[29][0],s2[29][1],s2[29][2],s3[29][1],c3[30][1]);
csa a3_30_0 (c2[30][0],c2[30][1],c2[30][2],s3[30][0],c3[31][0]);
csa a3_30_1 (s2[30][0],s2[30][1],s2[30][2],s3[30][1],c3[31][1]);
csa a3_31_0 (c2[31][0],c2[31][1],c2[31][2],s3[31][0],c3[32][0]);
csa a3_31_1 (s2[31][0],s2[31][1],s2[31][2],s3[31][1],c3[32][1]);
csa a3_32_0 (c2[32][0],c2[32][1],c2[32][2],s3[32][0],c3[33][0]);
csa a3_32_1 (s2[32][0],s2[32][1],s2[32][2],s3[32][1],c3[33][1]);
csa a3_33_0 (c2[33][0],c2[33][1],c2[33][2],s3[33][0],c3[34][0]);
csa a3_33_1 (s2[33][0],s2[33][1],s2[33][2],s3[33][1],c3[34][1]);
csa a3_34_0 (c2[34][0],c2[34][1],c2[34][2],s3[34][0],c3[35][0]);
csa a3_34_1 (s2[34][0],s2[34][1],s2[34][2],s3[34][1],c3[35][1]);
csa a3_35_0 (c2[35][0],c2[35][1],c2[35][2],s3[35][0],c3[36][0]);
csa a3_35_1 (s2[35][0],s2[35][1],s0[35][4],s3[35][1],c3[36][1]);
csa a3_36_0 (c2[36][0],c2[36][1],s2[36][0],s3[36][0],c3[37][0]);
csa a3_36_1 (s2[36][1],p[25][11],zero,s3[36][1],c3[37][1]);
csa a3_37_0 (c2[37][0],c2[37][1],s2[37][0],s3[37][0],c3[38][0]);
csa a3_38_0 (c2[38][0],c2[38][1],s2[38][0],s3[38][0],c3[39][0]);
csa a3_39_0 (c2[39][0],c2[39][1],s2[39][0],s3[39][0],c3[40][0]);
csa a3_40_0 (c2[40][0],c2[40][1],s2[40][0],s3[40][0],c3[41][0]);
csa a3_41_0 (c2[41][0],c2[41][1],s2[41][0],s3[41][0],c3[42][0]);
csa a3_42_0 (c2[42][0],s2[42][0],s1[42][1],s3[42][0],c3[43][0]);
csa a3_43_0 (c2[43][0],s2[43][0],s0[43][1],s3[43][0],c3[44][0]);
csa a3_44_0 (c2[44][0],s2[44][0],zero,s3[44][0],c3[45][0]);
csa a3_45_0 (c2[45][0],s2[45][0],zero,s3[45][0],c3[46][0]);
csa a3_46_0 (c2[46][0],s2[46][0],zero,s3[46][0],c3[47][0]);
csa a3_47_0 (c2[47][0],s2[47][0],zero,s3[47][0],c3[48][0]);
csa a3_48_0 (c2[48][0],s2[48][0],zero,s3[48][0],c3[49][0]);
csa a3_49_0 (c2[49][0],c1[49][0],zero,s3[49][0],c_overflow);

// level 4
wire [1:0] s4[0:49];
wire [1:0] c4[0:49];
csa a4_5_0 (c3[5][0],s3[5][0],zero,s4[5][0],c4[6][0]);
csa a4_6_0 (c3[6][0],s3[6][0],zero,s4[6][0],c4[7][0]);
csa a4_7_0 (c3[7][0],s3[7][0],zero,s4[7][0],c4[8][0]);
csa a4_8_0 (c3[8][0],s3[8][0],zero,s4[8][0],c4[9][0]);
csa a4_9_0 (c3[9][0],s3[9][0],zero,s4[9][0],c4[10][0]);
csa a4_10_0 (c3[10][0],s3[10][0],s2[10][1],s4[10][0],c4[11][0]);
csa a4_11_0 (c3[11][0],s3[11][0],s2[11][1],s4[11][0],c4[12][0]);
csa a4_12_0 (c3[12][0],s3[12][0],s2[12][1],s4[12][0],c4[13][0]);
csa a4_13_0 (c3[13][0],s3[13][0],s2[13][1],s4[13][0],c4[14][0]);
csa a4_14_0 (c3[14][0],s3[14][0],s3[14][1],s4[14][0],c4[15][0]);
csa a4_15_0 (c3[15][0],c3[15][1],s3[15][0],s4[15][0],c4[16][0]);
csa a4_16_0 (c3[16][0],c3[16][1],s3[16][0],s4[16][0],c4[17][0]);
csa a4_17_0 (c3[17][0],c3[17][1],s3[17][0],s4[17][0],c4[18][0]);
csa a4_18_0 (c3[18][0],c3[18][1],s3[18][0],s4[18][0],c4[19][0]);
csa a4_19_0 (c3[19][0],c3[19][1],s3[19][0],s4[19][0],c4[20][0]);
csa a4_20_0 (c3[20][0],c3[20][1],s3[20][0],s4[20][0],c4[21][0]);
csa a4_21_0 (c3[21][0],c3[21][1],s3[21][0],s4[21][0],c4[22][0]);
csa a4_21_1 (s3[21][1],s1[21][4],zero,s4[21][1],c4[22][1]);
csa a4_22_0 (c3[22][0],c3[22][1],s3[22][0],s4[22][0],c4[23][0]);
csa a4_22_1 (s3[22][1],s1[22][4],zero,s4[22][1],c4[23][1]);
csa a4_23_0 (c3[23][0],c3[23][1],s3[23][0],s4[23][0],c4[24][0]);
csa a4_23_1 (s3[23][1],s2[23][3],zero,s4[23][1],c4[24][1]);
csa a4_24_0 (c3[24][0],c3[24][1],s3[24][0],s4[24][0],c4[25][0]);
csa a4_24_1 (s3[24][1],s3[24][2],zero,s4[24][1],c4[25][1]);
csa a4_25_0 (c3[25][0],c3[25][1],c3[25][2],s4[25][0],c4[26][0]);
csa a4_25_1 (s3[25][0],s3[25][1],s3[25][2],s4[25][1],c4[26][1]);
csa a4_26_0 (c3[26][0],c3[26][1],c3[26][2],s4[26][0],c4[27][0]);
csa a4_26_1 (s3[26][0],s3[26][1],s3[26][2],s4[26][1],c4[27][1]);
csa a4_27_0 (c3[27][0],c3[27][1],c3[27][2],s4[27][0],c4[28][0]);
csa a4_27_1 (s3[27][0],s3[27][1],s3[27][2],s4[27][1],c4[28][1]);
csa a4_28_0 (c3[28][0],c3[28][1],c3[28][2],s4[28][0],c4[29][0]);
csa a4_28_1 (s3[28][0],s3[28][1],s3[28][2],s4[28][1],c4[29][1]);
csa a4_29_0 (c3[29][0],c3[29][1],c3[29][2],s4[29][0],c4[30][0]);
csa a4_29_1 (s3[29][0],s3[29][1],s1[29][4],s4[29][1],c4[30][1]);
csa a4_30_0 (c3[30][0],c3[30][1],s3[30][0],s4[30][0],c4[31][0]);
csa a4_30_1 (s3[30][1],s1[30][4],zero,s4[30][1],c4[31][1]);
csa a4_31_0 (c3[31][0],c3[31][1],s3[31][0],s4[31][0],c4[32][0]);
csa a4_32_0 (c3[32][0],c3[32][1],s3[32][0],s4[32][0],c4[33][0]);
csa a4_33_0 (c3[33][0],c3[33][1],s3[33][0],s4[33][0],c4[34][0]);
csa a4_34_0 (c3[34][0],c3[34][1],s3[34][0],s4[34][0],c4[35][0]);
csa a4_35_0 (c3[35][0],c3[35][1],s3[35][0],s4[35][0],c4[36][0]);
csa a4_36_0 (c3[36][0],c3[36][1],s3[36][0],s4[36][0],c4[37][0]);
csa a4_37_0 (c3[37][0],c3[37][1],s3[37][0],s4[37][0],c4[38][0]);
csa a4_38_0 (c3[38][0],s3[38][0],s2[38][1],s4[38][0],c4[39][0]);
csa a4_39_0 (c3[39][0],s3[39][0],s2[39][1],s4[39][0],c4[40][0]);
csa a4_40_0 (c3[40][0],s3[40][0],s2[40][1],s4[40][0],c4[41][0]);
csa a4_41_0 (c3[41][0],s3[41][0],s1[41][1],s4[41][0],c4[42][0]);
csa a4_42_0 (c3[42][0],s3[42][0],zero,s4[42][0],c4[43][0]);
csa a4_43_0 (c3[43][0],s3[43][0],zero,s4[43][0],c4[44][0]);
csa a4_44_0 (c3[44][0],s3[44][0],zero,s4[44][0],c4[45][0]);
csa a4_45_0 (c3[45][0],s3[45][0],zero,s4[45][0],c4[46][0]);
csa a4_46_0 (c3[46][0],s3[46][0],zero,s4[46][0],c4[47][0]);
csa a4_47_0 (c3[47][0],s3[47][0],zero,s4[47][0],c4[48][0]);
csa a4_48_0 (c3[48][0],s3[48][0],zero,s4[48][0],c4[49][0]);
csa a4_49_0 (c3[49][0],s3[49][0],zero,s4[49][0],c_overflow);

// level 5
wire [0:0] s5[0:49];
wire [0:0] c5[0:49];
csa a5_6_0 (c4[6][0],s4[6][0],zero,s5[6][0],c5[7][0]);
csa a5_7_0 (c4[7][0],s4[7][0],zero,s5[7][0],c5[8][0]);
csa a5_8_0 (c4[8][0],s4[8][0],zero,s5[8][0],c5[9][0]);
csa a5_9_0 (c4[9][0],s4[9][0],zero,s5[9][0],c5[10][0]);
csa a5_10_0 (c4[10][0],s4[10][0],zero,s5[10][0],c5[11][0]);
csa a5_11_0 (c4[11][0],s4[11][0],zero,s5[11][0],c5[12][0]);
csa a5_12_0 (c4[12][0],s4[12][0],zero,s5[12][0],c5[13][0]);
csa a5_13_0 (c4[13][0],s4[13][0],zero,s5[13][0],c5[14][0]);
csa a5_14_0 (c4[14][0],s4[14][0],zero,s5[14][0],c5[15][0]);
csa a5_15_0 (c4[15][0],s4[15][0],s3[15][1],s5[15][0],c5[16][0]);
csa a5_16_0 (c4[16][0],s4[16][0],s3[16][1],s5[16][0],c5[17][0]);
csa a5_17_0 (c4[17][0],s4[17][0],s3[17][1],s5[17][0],c5[18][0]);
csa a5_18_0 (c4[18][0],s4[18][0],s3[18][1],s5[18][0],c5[19][0]);
csa a5_19_0 (c4[19][0],s4[19][0],s3[19][1],s5[19][0],c5[20][0]);
csa a5_20_0 (c4[20][0],s4[20][0],s3[20][1],s5[20][0],c5[21][0]);
csa a5_21_0 (c4[21][0],s4[21][0],s4[21][1],s5[21][0],c5[22][0]);
csa a5_22_0 (c4[22][0],c4[22][1],s4[22][0],s5[22][0],c5[23][0]);
csa a5_23_0 (c4[23][0],c4[23][1],s4[23][0],s5[23][0],c5[24][0]);
csa a5_24_0 (c4[24][0],c4[24][1],s4[24][0],s5[24][0],c5[25][0]);
csa a5_25_0 (c4[25][0],c4[25][1],s4[25][0],s5[25][0],c5[26][0]);
csa a5_26_0 (c4[26][0],c4[26][1],s4[26][0],s5[26][0],c5[27][0]);
csa a5_27_0 (c4[27][0],c4[27][1],s4[27][0],s5[27][0],c5[28][0]);
csa a5_28_0 (c4[28][0],c4[28][1],s4[28][0],s5[28][0],c5[29][0]);
csa a5_29_0 (c4[29][0],c4[29][1],s4[29][0],s5[29][0],c5[30][0]);
csa a5_30_0 (c4[30][0],c4[30][1],s4[30][0],s5[30][0],c5[31][0]);
csa a5_31_0 (c4[31][0],c4[31][1],s4[31][0],s5[31][0],c5[32][0]);
csa a5_32_0 (c4[32][0],s4[32][0],s3[32][1],s5[32][0],c5[33][0]);
csa a5_33_0 (c4[33][0],s4[33][0],s3[33][1],s5[33][0],c5[34][0]);
csa a5_34_0 (c4[34][0],s4[34][0],s3[34][1],s5[34][0],c5[35][0]);
csa a5_35_0 (c4[35][0],s4[35][0],s3[35][1],s5[35][0],c5[36][0]);
csa a5_36_0 (c4[36][0],s4[36][0],s3[36][1],s5[36][0],c5[37][0]);
csa a5_37_0 (c4[37][0],s4[37][0],s2[37][1],s5[37][0],c5[38][0]);
csa a5_38_0 (c4[38][0],s4[38][0],zero,s5[38][0],c5[39][0]);
csa a5_39_0 (c4[39][0],s4[39][0],zero,s5[39][0],c5[40][0]);
csa a5_40_0 (c4[40][0],s4[40][0],zero,s5[40][0],c5[41][0]);
csa a5_41_0 (c4[41][0],s4[41][0],zero,s5[41][0],c5[42][0]);
csa a5_42_0 (c4[42][0],s4[42][0],zero,s5[42][0],c5[43][0]);
csa a5_43_0 (c4[43][0],s4[43][0],zero,s5[43][0],c5[44][0]);
csa a5_44_0 (c4[44][0],s4[44][0],zero,s5[44][0],c5[45][0]);
csa a5_45_0 (c4[45][0],s4[45][0],zero,s5[45][0],c5[46][0]);
csa a5_46_0 (c4[46][0],s4[46][0],zero,s5[46][0],c5[47][0]);
csa a5_47_0 (c4[47][0],s4[47][0],zero,s5[47][0],c5[48][0]);
csa a5_48_0 (c4[48][0],s4[48][0],zero,s5[48][0],c5[49][0]);
csa a5_49_0 (c4[49][0],s4[49][0],zero,s5[49][0],c_overflow);

// level 6
wire [0:0] s6[0:49];
wire [0:0] c6[0:49];
csa a6_7_0 (c5[7][0],s5[7][0],zero,s6[7][0],c6[8][0]);
csa a6_8_0 (c5[8][0],s5[8][0],zero,s6[8][0],c6[9][0]);
csa a6_9_0 (c5[9][0],s5[9][0],zero,s6[9][0],c6[10][0]);
csa a6_10_0 (c5[10][0],s5[10][0],zero,s6[10][0],c6[11][0]);
csa a6_11_0 (c5[11][0],s5[11][0],zero,s6[11][0],c6[12][0]);
csa a6_12_0 (c5[12][0],s5[12][0],zero,s6[12][0],c6[13][0]);
csa a6_13_0 (c5[13][0],s5[13][0],zero,s6[13][0],c6[14][0]);
csa a6_14_0 (c5[14][0],s5[14][0],zero,s6[14][0],c6[15][0]);
csa a6_15_0 (c5[15][0],s5[15][0],zero,s6[15][0],c6[16][0]);
csa a6_16_0 (c5[16][0],s5[16][0],zero,s6[16][0],c6[17][0]);
csa a6_17_0 (c5[17][0],s5[17][0],zero,s6[17][0],c6[18][0]);
csa a6_18_0 (c5[18][0],s5[18][0],zero,s6[18][0],c6[19][0]);
csa a6_19_0 (c5[19][0],s5[19][0],zero,s6[19][0],c6[20][0]);
csa a6_20_0 (c5[20][0],s5[20][0],zero,s6[20][0],c6[21][0]);
csa a6_21_0 (c5[21][0],s5[21][0],zero,s6[21][0],c6[22][0]);
csa a6_22_0 (c5[22][0],s5[22][0],s4[22][1],s6[22][0],c6[23][0]);
csa a6_23_0 (c5[23][0],s5[23][0],s4[23][1],s6[23][0],c6[24][0]);
csa a6_24_0 (c5[24][0],s5[24][0],s4[24][1],s6[24][0],c6[25][0]);
csa a6_25_0 (c5[25][0],s5[25][0],s4[25][1],s6[25][0],c6[26][0]);
csa a6_26_0 (c5[26][0],s5[26][0],s4[26][1],s6[26][0],c6[27][0]);
csa a6_27_0 (c5[27][0],s5[27][0],s4[27][1],s6[27][0],c6[28][0]);
csa a6_28_0 (c5[28][0],s5[28][0],s4[28][1],s6[28][0],c6[29][0]);
csa a6_29_0 (c5[29][0],s5[29][0],s4[29][1],s6[29][0],c6[30][0]);
csa a6_30_0 (c5[30][0],s5[30][0],s4[30][1],s6[30][0],c6[31][0]);
csa a6_31_0 (c5[31][0],s5[31][0],s3[31][1],s6[31][0],c6[32][0]);
csa a6_32_0 (c5[32][0],s5[32][0],zero,s6[32][0],c6[33][0]);
csa a6_33_0 (c5[33][0],s5[33][0],zero,s6[33][0],c6[34][0]);
csa a6_34_0 (c5[34][0],s5[34][0],zero,s6[34][0],c6[35][0]);
csa a6_35_0 (c5[35][0],s5[35][0],zero,s6[35][0],c6[36][0]);
csa a6_36_0 (c5[36][0],s5[36][0],zero,s6[36][0],c6[37][0]);
csa a6_37_0 (c5[37][0],s5[37][0],zero,s6[37][0],c6[38][0]);
csa a6_38_0 (c5[38][0],s5[38][0],zero,s6[38][0],c6[39][0]);
csa a6_39_0 (c5[39][0],s5[39][0],zero,s6[39][0],c6[40][0]);
csa a6_40_0 (c5[40][0],s5[40][0],zero,s6[40][0],c6[41][0]);
csa a6_41_0 (c5[41][0],s5[41][0],zero,s6[41][0],c6[42][0]);
csa a6_42_0 (c5[42][0],s5[42][0],zero,s6[42][0],c6[43][0]);
csa a6_43_0 (c5[43][0],s5[43][0],zero,s6[43][0],c6[44][0]);
csa a6_44_0 (c5[44][0],s5[44][0],zero,s6[44][0],c6[45][0]);
csa a6_45_0 (c5[45][0],s5[45][0],zero,s6[45][0],c6[46][0]);
csa a6_46_0 (c5[46][0],s5[46][0],zero,s6[46][0],c6[47][0]);
csa a6_47_0 (c5[47][0],s5[47][0],zero,s6[47][0],c6[48][0]);
csa a6_48_0 (c5[48][0],s5[48][0],zero,s6[48][0],c6[49][0]);
csa a6_49_0 (c5[49][0],s5[49][0],zero,s6[49][0],c_overflow);

// final assignment to x, y, z
assign z[0] = p[0][0];
assign z[1] = s0[1][0];
assign z[2] = s1[2][0];
assign z[3] = s2[3][0];
assign z[4] = s3[4][0];
assign z[5] = s4[5][0];
assign z[6] = s5[6][0];
assign z[7] = s6[7][0];
assign x[8] = c6[8][0];
assign y[8] = s6[8][0];
assign x[9] = c6[9][0];
assign y[9] = s6[9][0];
assign x[10] = c6[10][0];
assign y[10] = s6[10][0];
assign x[11] = c6[11][0];
assign y[11] = s6[11][0];
assign x[12] = c6[12][0];
assign y[12] = s6[12][0];
assign x[13] = c6[13][0];
assign y[13] = s6[13][0];
assign x[14] = c6[14][0];
assign y[14] = s6[14][0];
assign x[15] = c6[15][0];
assign y[15] = s6[15][0];
assign x[16] = c6[16][0];
assign y[16] = s6[16][0];
assign x[17] = c6[17][0];
assign y[17] = s6[17][0];
assign x[18] = c6[18][0];
assign y[18] = s6[18][0];
assign x[19] = c6[19][0];
assign y[19] = s6[19][0];
assign x[20] = c6[20][0];
assign y[20] = s6[20][0];
assign x[21] = c6[21][0];
assign y[21] = s6[21][0];
assign x[22] = c6[22][0];
assign y[22] = s6[22][0];
assign x[23] = c6[23][0];
assign y[23] = s6[23][0];
assign x[24] = c6[24][0];
assign y[24] = s6[24][0];
assign x[25] = c6[25][0];
assign y[25] = s6[25][0];
assign x[26] = c6[26][0];
assign y[26] = s6[26][0];
assign x[27] = c6[27][0];
assign y[27] = s6[27][0];
assign x[28] = c6[28][0];
assign y[28] = s6[28][0];
assign x[29] = c6[29][0];
assign y[29] = s6[29][0];
assign x[30] = c6[30][0];
assign y[30] = s6[30][0];
assign x[31] = c6[31][0];
assign y[31] = s6[31][0];
assign x[32] = c6[32][0];
assign y[32] = s6[32][0];
assign x[33] = c6[33][0];
assign y[33] = s6[33][0];
assign x[34] = c6[34][0];
assign y[34] = s6[34][0];
assign x[35] = c6[35][0];
assign y[35] = s6[35][0];
assign x[36] = c6[36][0];
assign y[36] = s6[36][0];
assign x[37] = c6[37][0];
assign y[37] = s6[37][0];
assign x[38] = c6[38][0];
assign y[38] = s6[38][0];
assign x[39] = c6[39][0];
assign y[39] = s6[39][0];
assign x[40] = c6[40][0];
assign y[40] = s6[40][0];
assign x[41] = c6[41][0];
assign y[41] = s6[41][0];
assign x[42] = c6[42][0];
assign y[42] = s6[42][0];
assign x[43] = c6[43][0];
assign y[43] = s6[43][0];
assign x[44] = c6[44][0];
assign y[44] = s6[44][0];
assign x[45] = c6[45][0];
assign y[45] = s6[45][0];
assign x[46] = c6[46][0];
assign y[46] = s6[46][0];
assign x[47] = c6[47][0];
assign y[47] = s6[47][0];
assign x[48] = c6[48][0];
assign y[48] = s6[48][0];
assign x[49] = c6[49][0];
assign y[49] = s6[49][0];

endmodule
